magic
tech scmos
timestamp 1701337605
<< polysilicon >>
rect -20 63 -18 70
rect -100 61 -18 63
rect -100 58 -98 61
rect -20 58 -18 61
rect 11 63 13 70
rect 11 61 94 63
rect 11 58 13 61
rect 92 58 94 61
rect -110 2 -108 6
rect 11 2 13 5
rect -110 0 13 2
<< polycontact >>
rect -21 70 -17 74
rect 10 70 14 74
<< metal1 >>
rect -21 74 -17 78
rect 10 74 14 78
rect -6 64 0 67
rect 19 39 25 43
rect -6 0 0 4
rect -140 -15 -135 -10
rect -85 -15 -80 -10
rect 74 -15 79 -10
rect 129 -15 134 -10
<< m2contact >>
rect -36 27 -31 32
rect -12 27 -7 32
rect 25 27 30 32
rect 80 27 85 32
rect -140 15 -135 20
rect -85 15 -80 20
rect 15 18 20 23
rect 74 15 79 20
rect 129 15 134 20
rect -140 -10 -135 -5
rect -85 -10 -80 -5
rect 74 -10 79 -5
rect 129 -10 134 -5
<< metal2 >>
rect -7 27 25 32
rect 30 27 80 32
rect -36 23 -31 27
rect -140 -5 -135 15
rect -36 18 15 23
rect -85 -5 -80 15
rect 74 -5 79 15
rect 129 -5 134 15
use NOT  NOT_0
timestamp 1701333315
transform 1 0 36 0 1 2
box -36 -2 -11 65
use NOT  NOT_1
timestamp 1701333315
transform 1 0 5 0 1 2
box -36 -2 -11 65
use AND  AND_0
timestamp 1701179155
transform 1 0 -39 0 1 0
box 64 0 119 67
use AND  AND_1
timestamp 1701179155
transform 1 0 16 0 1 0
box 64 0 119 67
use AND  AND_2
timestamp 1701179155
transform -1 0 33 0 1 0
box 64 0 119 67
use AND  AND_3
timestamp 1701179155
transform -1 0 -22 0 1 0
box 64 0 119 67
<< labels >>
rlabel metal1 -3 65 -3 65 5 vdd
rlabel metal1 -3 1 -3 1 1 gnd
rlabel metal1 -19 76 -19 76 5 S0
rlabel metal1 12 76 12 76 5 S1
rlabel metal1 76 -13 76 -13 1 R0
rlabel metal1 131 -13 131 -13 8 R2
rlabel metal1 -83 -13 -83 -13 1 R1
rlabel metal1 -138 -13 -138 -13 2 R3
<< end >>
