*CMOS Half Adder

.include TSMC_180nm.txt
.param supply=1.5
.option scale=0.09u

V1 vdd gnd supply

M1000 NAND_0/out B NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1001 NAND_0/out A vdd vdd CMOSP w=4 l=2
+  ad=32 pd=24 as=176 ps=144
M1002 vdd B NAND_0/out vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 NAND_0/a_n7_n34# A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=152 ps=124
M1004 Sum A XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1005 XOR_0/a_123_36# A vdd vdd CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1006 Sum B XOR_0/a_141_74# vdd CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1007 XOR_0/a_141_36# B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 gnd XOR_0/a_184_44# XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1009 XOR_0/a_141_74# XOR_0/a_123_36# vdd vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 vdd XOR_0/a_184_44# XOR_0/a_177_74# vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1011 XOR_0/a_177_36# XOR_0/a_123_36# Sum Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 XOR_0/a_177_74# A Sum vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 gnd B XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1014 vdd B XOR_0/a_184_44# vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1015 XOR_0/a_123_36# A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1016 Cout NAND_0/out vdd vdd CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1017 Cout NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
C0 vdd XOR_0/a_123_36# 0.09fF
C1 A NAND_0/out 0.14fF
C2 Sum XOR_0/a_141_36# 0.03fF
C3 vdd B 0.70fF
C4 Sum B 0.11fF
C5 vdd vdd 0.22fF
C6 vdd B 0.29fF
C7 NAND_0/out Cout 0.05fF
C8 vdd XOR_0/a_177_74# 0.01fF
C9 vdd vdd 0.14fF
C10 Sum XOR_0/a_177_74# 0.03fF
C11 Sum XOR_0/a_177_36# 0.03fF
C12 A vdd 0.13fF
C13 A Sum 0.23fF
C14 vdd XOR_0/a_141_74# 0.01fF
C15 vdd A 0.06fF
C16 XOR_0/a_141_74# Sum 0.03fF
C17 XOR_0/a_123_36# B 0.10fF
C18 vdd XOR_0/a_123_36# 0.06fF
C19 vdd Cout 0.03fF
C20 vdd B 0.32fF
C21 vdd XOR_0/a_184_44# 0.09fF
C22 XOR_0/a_184_44# Sum 0.13fF
C23 gnd XOR_0/a_123_36# 0.14fF
C24 gnd XOR_0/a_141_36# 0.02fF
C25 A XOR_0/a_123_36# 0.26fF
C26 A XOR_0/a_141_36# 0.03fF
C27 vdd XOR_0/a_177_74# 0.02fF
C28 A B 0.59fF
C29 vdd NAND_0/out 0.09fF
C30 gnd XOR_0/a_177_36# 0.02fF
C31 vdd XOR_0/a_141_74# 0.02fF
C32 vdd Cout 0.03fF
C33 A gnd 0.03fF
C34 vdd Sum 0.06fF
C35 XOR_0/a_184_44# B 0.06fF
C36 gnd Cout 0.07fF
C37 vdd XOR_0/a_184_44# 0.06fF
C38 A Cout 0.10fF
C39 NAND_0/out B 0.20fF
C40 vdd NAND_0/out 0.06fF
C41 gnd XOR_0/a_184_44# 0.11fF
C42 A XOR_0/a_184_44# 0.00fF
C43 NAND_0/out gnd 0.04fF
C44 Cout Gnd 0.13fF
C45 B Gnd 1.07fF
C46 XOR_0/a_177_36# Gnd 0.01fF
C47 XOR_0/a_141_36# Gnd 0.01fF
C48 Sum Gnd 0.34fF
C49 XOR_0/a_184_44# Gnd 0.34fF
C50 XOR_0/a_123_36# Gnd 0.80fF
C51 vdd Gnd 2.10fF
C52 gnd Gnd 0.52fF
C53 NAND_0/out Gnd 0.43fF
C54 vdd Gnd 0.28fF
C55 A Gnd 2.28fF
C56 vdd Gnd 1.11fF

Vin1 A GND pulse(0 supply 0 0.5p 0.5p 0.1u 0.2u)
Vin2 B GND pulse(0 supply 0.15u 0.5p 0.5p 0.1u 0.2u)

.control
tran 1p 0.4u
plot v(A) v(B)+3 V(Sum)+6 V(Cout)+9
.endc
.end