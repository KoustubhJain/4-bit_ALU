*Four Bit CMOS ALU

.include TSMC_180nm.txt
.param supply=1.5
.option scale=0.09u

V1 vdd gnd supply

M1000 gnd ALU_1b_0/NOR_2/B ALU_1b_0/NOT_4/in Gnd CMOSN w=4 l=2
+  ad=11824 pd=9848 as=24 ps=20
M1001 ALU_1b_0/NOT_4/in ALU_1b_0/NOR_2/B ALU_1b_0/NOR_2/a_n14_7# ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1002 ALU_1b_0/NOR_2/a_n14_7# ALU_1b_0/NOR_2/A vdd ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=13764 ps=11524
M1003 ALU_1b_0/NOT_4/in ALU_1b_0/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 ALU_1b_0/NOR_4/B ALU_1b_0/NOT_5/in vdd ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1005 ALU_1b_0/NOR_4/B ALU_1b_0/NOT_5/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1006 ALU_1b_2/C0 ALU_1b_0/NOT_6/in vdd ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1007 ALU_1b_2/C0 ALU_1b_0/NOT_6/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1008 gnd ALU_1b_0/NOR_3/B ALU_1b_0/NOT_5/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1009 ALU_1b_0/NOT_5/in ALU_1b_0/NOR_3/B ALU_1b_0/NOR_3/a_n14_7# ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1010 ALU_1b_0/NOR_3/a_n14_7# ALU_1b_0/NOR_3/A vdd ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 ALU_1b_0/NOT_5/in ALU_1b_0/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 gnd ALU_1b_0/NOR_4/B ALU_1b_0/NOT_6/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1013 ALU_1b_0/NOT_6/in ALU_1b_0/NOR_4/B ALU_1b_0/NOR_4/a_n14_7# ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1014 ALU_1b_0/NOR_4/a_n14_7# ALU_1b_0/NOR_4/A vdd ALU_1b_0/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1015 ALU_1b_0/NOT_6/in ALU_1b_0/NOR_4/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1016 ALU_1b_0/AND_0/a_78_51# A0 ALU_1b_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1017 ALU_1b_0/AND_0/out ALU_1b_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1018 vdd A0 ALU_1b_0/AND_0/a_78_51# ALU_1b_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1019 ALU_1b_0/AND_0/a_78_51# ALU_1b_0/AND_2/B vdd ALU_1b_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1020 ALU_1b_0/AND_0/a_78_8# ALU_1b_0/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1021 ALU_1b_0/AND_0/out ALU_1b_0/AND_0/a_78_51# vdd ALU_1b_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1022 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1023 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/full_adder_0/half_adder_1/A vdd ALU_1b_0/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1024 vdd ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1025 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/a_n7_n34# ALU_1b_0/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1026 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1027 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_0/half_adder_1/A vdd ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1028 ALU_1b_0/AND_16/A ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1029 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_0/AND_1/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1030 gnd ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1031 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1032 vdd ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1033 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/AND_16/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 gnd ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1036 vdd ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1037 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1038 ALU_1b_0/full_adder_0/NOR_0/A ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out vdd ALU_1b_0/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1039 ALU_1b_0/full_adder_0/NOR_0/A ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1040 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1041 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/AND_0/out vdd ALU_1b_0/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1042 vdd ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_0/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1045 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_0/out vdd ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1046 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1047 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# ALU_1b_0/AND_2/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1048 gnd ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1049 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1050 vdd ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1051 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_0/full_adder_0/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1052 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1053 gnd ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1054 vdd ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1055 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1056 ALU_1b_0/full_adder_0/NOR_0/B ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out vdd ALU_1b_0/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1057 ALU_1b_0/full_adder_0/NOR_0/B ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1058 gnd ALU_1b_0/full_adder_0/NOR_0/B ALU_1b_0/full_adder_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1059 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/full_adder_0/NOR_0/B ALU_1b_0/full_adder_0/NOR_0/a_n14_7# ALU_1b_0/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1060 ALU_1b_0/full_adder_0/NOR_0/a_n14_7# ALU_1b_0/full_adder_0/NOR_0/A vdd ALU_1b_0/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/full_adder_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 ALU_1b_0/AND_17/A ALU_1b_0/full_adder_0/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1063 ALU_1b_0/AND_17/A ALU_1b_0/full_adder_0/NOR_0/out vdd ALU_1b_0/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1064 ALU_1b_0/AND_1/a_78_51# ALU_1b_0/AND_2/B ALU_1b_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1065 ALU_1b_0/AND_1/out ALU_1b_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1066 vdd ALU_1b_0/AND_2/B ALU_1b_0/AND_1/a_78_51# ALU_1b_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1067 ALU_1b_0/AND_1/a_78_51# Cin vdd ALU_1b_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 ALU_1b_0/AND_1/a_78_8# Cin gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1069 ALU_1b_0/AND_1/out ALU_1b_0/AND_1/a_78_51# vdd ALU_1b_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1070 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1071 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/full_adder_1/half_adder_1/A vdd ALU_1b_0/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1072 vdd ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1073 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/a_n7_n34# ALU_1b_0/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1075 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_1/half_adder_1/A vdd ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1076 ALU_1b_0/NOT_1/in ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1077 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_0/AND_5/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1078 gnd ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1079 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 vdd ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1081 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/NOT_1/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1083 gnd ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1084 vdd ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1085 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1086 ALU_1b_0/full_adder_1/NOR_0/A ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out vdd ALU_1b_0/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1087 ALU_1b_0/full_adder_1/NOR_0/A ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1088 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1089 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/AND_3/out vdd ALU_1b_0/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1090 vdd ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1091 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_0/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1092 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1093 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_3/out vdd ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1094 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1095 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_0/AND_4/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 gnd ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1097 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1098 vdd ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1099 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_0/full_adder_1/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 gnd ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1102 vdd ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1103 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1104 ALU_1b_0/full_adder_1/NOR_0/B ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out vdd ALU_1b_0/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1105 ALU_1b_0/full_adder_1/NOR_0/B ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1106 gnd ALU_1b_0/full_adder_1/NOR_0/B ALU_1b_0/full_adder_1/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1107 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/full_adder_1/NOR_0/B ALU_1b_0/full_adder_1/NOR_0/a_n14_7# ALU_1b_0/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1108 ALU_1b_0/full_adder_1/NOR_0/a_n14_7# ALU_1b_0/full_adder_1/NOR_0/A vdd ALU_1b_0/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/full_adder_1/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 ALU_1b_0/AND_18/A ALU_1b_0/full_adder_1/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1111 ALU_1b_0/AND_18/A ALU_1b_0/full_adder_1/NOR_0/out vdd ALU_1b_0/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1112 ALU_1b_0/AND_2/a_78_51# ALU_1b_0/AND_2/B ALU_1b_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1113 ALU_1b_0/AND_2/out ALU_1b_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1114 vdd ALU_1b_0/AND_2/B ALU_1b_0/AND_2/a_78_51# ALU_1b_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1115 ALU_1b_0/AND_2/a_78_51# B0 vdd ALU_1b_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1116 ALU_1b_0/AND_2/a_78_8# B0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1117 ALU_1b_0/AND_2/out ALU_1b_0/AND_2/a_78_51# vdd ALU_1b_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1118 ALU_1b_0/AND_3/a_78_51# ALU_1b_0/AND_5/B ALU_1b_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1119 ALU_1b_0/AND_3/out ALU_1b_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1120 vdd ALU_1b_0/AND_5/B ALU_1b_0/AND_3/a_78_51# ALU_1b_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1121 ALU_1b_0/AND_3/a_78_51# ALU_1b_0/AND_3/A vdd ALU_1b_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1122 ALU_1b_0/AND_3/a_78_8# ALU_1b_0/AND_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 ALU_1b_0/AND_3/out ALU_1b_0/AND_3/a_78_51# vdd ALU_1b_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1124 ALU_1b_0/AND_5/a_78_51# ALU_1b_0/AND_5/B ALU_1b_0/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1125 ALU_1b_0/AND_5/out ALU_1b_0/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1126 vdd ALU_1b_0/AND_5/B ALU_1b_0/AND_5/a_78_51# ALU_1b_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1127 ALU_1b_0/AND_5/a_78_51# Cin vdd ALU_1b_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 ALU_1b_0/AND_5/a_78_8# Cin gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 ALU_1b_0/AND_5/out ALU_1b_0/AND_5/a_78_51# vdd ALU_1b_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1130 ALU_1b_0/AND_4/a_78_51# ALU_1b_0/AND_5/B ALU_1b_0/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1131 ALU_1b_0/AND_4/out ALU_1b_0/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1132 vdd ALU_1b_0/AND_5/B ALU_1b_0/AND_4/a_78_51# ALU_1b_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1133 ALU_1b_0/AND_4/a_78_51# B0 vdd ALU_1b_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 ALU_1b_0/AND_4/a_78_8# B0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1135 ALU_1b_0/AND_4/out ALU_1b_0/AND_4/a_78_51# vdd ALU_1b_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1136 ALU_1b_0/AND_10/a_78_51# ALU_1b_0/AND_10/B ALU_1b_0/AND_10/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1137 ALU_1b_0/NOR_1/A ALU_1b_0/AND_10/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1138 vdd ALU_1b_0/AND_10/B ALU_1b_0/AND_10/a_78_51# ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1139 ALU_1b_0/AND_10/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 ALU_1b_0/AND_10/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 ALU_1b_0/NOR_1/A ALU_1b_0/AND_10/a_78_51# vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1142 ALU_1b_0/AND_11/a_78_51# ALU_1b_0/AND_11/B ALU_1b_0/AND_11/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1143 ALU_1b_0/NOR_4/A ALU_1b_0/AND_11/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1144 vdd ALU_1b_0/AND_11/B ALU_1b_0/AND_11/a_78_51# ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1145 ALU_1b_0/AND_11/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1146 ALU_1b_0/AND_11/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 ALU_1b_0/NOR_4/A ALU_1b_0/AND_11/a_78_51# vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1148 ALU_1b_0/AND_6/a_78_51# A0 ALU_1b_0/AND_6/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1149 ALU_1b_0/AND_6/out ALU_1b_0/AND_6/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1150 vdd A0 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1151 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 ALU_1b_0/AND_6/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 ALU_1b_0/AND_6/out ALU_1b_0/AND_6/a_78_51# vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1154 ALU_1b_0/AND_7/a_78_51# B0 ALU_1b_0/AND_7/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1155 ALU_1b_0/AND_7/out ALU_1b_0/AND_7/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1156 vdd B0 ALU_1b_0/AND_7/a_78_51# ALU_1b_0/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1157 ALU_1b_0/AND_7/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1158 ALU_1b_0/AND_7/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 ALU_1b_0/AND_7/out ALU_1b_0/AND_7/a_78_51# vdd ALU_1b_0/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1160 ALU_1b_0/AND_12/a_78_51# A0 ALU_1b_0/AND_12/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1161 ALU_1b_0/AND_14/B ALU_1b_0/AND_12/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1162 vdd A0 ALU_1b_0/AND_12/a_78_51# ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1163 ALU_1b_0/AND_12/a_78_51# ALU_1b_0/AND_15/A vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1164 ALU_1b_0/AND_12/a_78_8# ALU_1b_0/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 ALU_1b_0/AND_14/B ALU_1b_0/AND_12/a_78_51# vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1166 ALU_1b_0/AND_8/a_78_51# C0 ALU_1b_0/AND_8/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1167 ALU_1b_0/AND_8/out ALU_1b_0/AND_8/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1168 vdd C0 ALU_1b_0/AND_8/a_78_51# ALU_1b_0/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1169 ALU_1b_0/AND_8/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 ALU_1b_0/AND_8/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1171 ALU_1b_0/AND_8/out ALU_1b_0/AND_8/a_78_51# vdd ALU_1b_0/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1172 ALU_1b_0/AND_13/a_78_51# B0 ALU_1b_0/AND_13/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1173 ALU_1b_0/AND_14/A ALU_1b_0/AND_13/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1174 vdd B0 ALU_1b_0/AND_13/a_78_51# ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1175 ALU_1b_0/AND_13/a_78_51# ALU_1b_0/AND_15/A vdd ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 ALU_1b_0/AND_13/a_78_8# ALU_1b_0/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 ALU_1b_0/AND_14/A ALU_1b_0/AND_13/a_78_51# vdd ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1178 ALU_1b_0/AND_9/a_78_51# C1 ALU_1b_0/AND_9/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1179 ALU_1b_0/AND_9/out ALU_1b_0/AND_9/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1180 vdd C1 ALU_1b_0/AND_9/a_78_51# ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1181 ALU_1b_0/AND_9/a_78_51# ALU_1b_0/AND_9/A vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 ALU_1b_0/AND_9/a_78_8# ALU_1b_0/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 ALU_1b_0/AND_9/out ALU_1b_0/AND_9/a_78_51# vdd ALU_1b_0/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1184 ALU_1b_0/AND_14/a_78_51# ALU_1b_0/AND_14/B ALU_1b_0/AND_14/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1185 ALU_1b_0/AND_15/B ALU_1b_0/AND_14/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1186 vdd ALU_1b_0/AND_14/B ALU_1b_0/AND_14/a_78_51# ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1187 ALU_1b_0/AND_14/a_78_51# ALU_1b_0/AND_14/A vdd ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 ALU_1b_0/AND_14/a_78_8# ALU_1b_0/AND_14/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 ALU_1b_0/AND_15/B ALU_1b_0/AND_14/a_78_51# vdd ALU_1b_0/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1190 ALU_1b_0/AND_15/a_78_51# ALU_1b_0/AND_15/B ALU_1b_0/AND_15/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1191 ALU_1b_0/NOR_1/B ALU_1b_0/AND_15/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1192 vdd ALU_1b_0/AND_15/B ALU_1b_0/AND_15/a_78_51# ALU_1b_0/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1193 ALU_1b_0/AND_15/a_78_51# ALU_1b_0/AND_15/A vdd ALU_1b_0/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 ALU_1b_0/AND_15/a_78_8# ALU_1b_0/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 ALU_1b_0/NOR_1/B ALU_1b_0/AND_15/a_78_51# vdd ALU_1b_0/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1196 ALU_1b_0/AND_16/a_78_51# ALU_1b_0/AND_2/B ALU_1b_0/AND_16/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1197 ALU_1b_0/NOR_0/B ALU_1b_0/AND_16/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1198 vdd ALU_1b_0/AND_2/B ALU_1b_0/AND_16/a_78_51# ALU_1b_0/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1199 ALU_1b_0/AND_16/a_78_51# ALU_1b_0/AND_16/A vdd ALU_1b_0/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 ALU_1b_0/AND_16/a_78_8# ALU_1b_0/AND_16/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1201 ALU_1b_0/NOR_0/B ALU_1b_0/AND_16/a_78_51# vdd ALU_1b_0/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1202 ALU_1b_0/AND_17/a_78_51# ALU_1b_0/AND_2/B ALU_1b_0/AND_17/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1203 ALU_1b_0/NOR_3/B ALU_1b_0/AND_17/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1204 vdd ALU_1b_0/AND_2/B ALU_1b_0/AND_17/a_78_51# ALU_1b_0/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1205 ALU_1b_0/AND_17/a_78_51# ALU_1b_0/AND_17/A vdd ALU_1b_0/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 ALU_1b_0/AND_17/a_78_8# ALU_1b_0/AND_17/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 ALU_1b_0/NOR_3/B ALU_1b_0/AND_17/a_78_51# vdd ALU_1b_0/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1208 ALU_1b_0/AND_19/a_78_51# ALU_1b_0/AND_5/B ALU_1b_0/AND_19/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1209 ALU_1b_0/NOR_0/A ALU_1b_0/AND_19/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1210 vdd ALU_1b_0/AND_5/B ALU_1b_0/AND_19/a_78_51# ALU_1b_0/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1211 ALU_1b_0/AND_19/a_78_51# ALU_1b_0/AND_19/A vdd ALU_1b_0/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 ALU_1b_0/AND_19/a_78_8# ALU_1b_0/AND_19/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 ALU_1b_0/NOR_0/A ALU_1b_0/AND_19/a_78_51# vdd ALU_1b_0/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1214 ALU_1b_0/AND_18/a_78_51# ALU_1b_0/AND_5/B ALU_1b_0/AND_18/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1215 ALU_1b_0/NOR_3/A ALU_1b_0/AND_18/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1216 vdd ALU_1b_0/AND_5/B ALU_1b_0/AND_18/a_78_51# ALU_1b_0/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1217 ALU_1b_0/AND_18/a_78_51# ALU_1b_0/AND_18/A vdd ALU_1b_0/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 ALU_1b_0/AND_18/a_78_8# ALU_1b_0/AND_18/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1219 ALU_1b_0/NOR_3/A ALU_1b_0/AND_18/a_78_51# vdd ALU_1b_0/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1220 gnd ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_2/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1221 ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_2/a_n14_7# ALU_1b_0/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1222 ALU_1b_0/comparator_0/NOR_2/a_n14_7# ALU_1b_0/comparator_0/NOR_2/A vdd ALU_1b_0/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/comparator_0/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 gnd ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/NOR_3/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1225 ALU_1b_0/comparator_0/NOR_3/out ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/NOR_3/a_n14_7# ALU_1b_0/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1226 ALU_1b_0/comparator_0/NOR_3/a_n14_7# ALU_1b_0/comparator_0/NOR_3/A vdd ALU_1b_0/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 ALU_1b_0/comparator_0/NOR_3/out ALU_1b_0/comparator_0/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 ALU_1b_0/comparator_0/AND_0/a_78_51# ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1229 ALU_1b_0/comparator_0/NOR_0/A ALU_1b_0/comparator_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1230 vdd ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_0/a_78_51# ALU_1b_0/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1231 ALU_1b_0/comparator_0/AND_0/a_78_51# ALU_1b_0/AND_6/out vdd ALU_1b_0/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 ALU_1b_0/comparator_0/AND_0/a_78_8# ALU_1b_0/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1233 ALU_1b_0/comparator_0/NOR_0/A ALU_1b_0/comparator_0/AND_0/a_78_51# vdd ALU_1b_0/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1234 ALU_1b_0/comparator_0/AND_1/a_78_51# ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1235 ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1236 vdd ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/AND_1/a_78_51# ALU_1b_0/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1237 ALU_1b_0/comparator_0/AND_1/a_78_51# ALU_1b_0/AND_6/out vdd ALU_1b_0/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 ALU_1b_0/comparator_0/AND_1/a_78_8# ALU_1b_0/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/AND_1/a_78_51# vdd ALU_1b_0/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1240 ALU_1b_0/comparator_0/AND_2/a_78_51# ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1241 ALU_1b_0/comparator_0/NOR_1/A ALU_1b_0/comparator_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1242 vdd ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_2/a_78_51# ALU_1b_0/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1243 ALU_1b_0/comparator_0/AND_2/a_78_51# ALU_1b_0/AND_9/out vdd ALU_1b_0/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1244 ALU_1b_0/comparator_0/AND_2/a_78_8# ALU_1b_0/AND_9/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1245 ALU_1b_0/comparator_0/NOR_1/A ALU_1b_0/comparator_0/AND_2/a_78_51# vdd ALU_1b_0/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1246 ALU_1b_0/comparator_0/AND_3/a_78_51# ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1247 ALU_1b_0/comparator_0/NOR_2/A ALU_1b_0/comparator_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1248 vdd ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_3/a_78_51# ALU_1b_0/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1249 ALU_1b_0/comparator_0/AND_3/a_78_51# ALU_1b_0/AND_8/out vdd ALU_1b_0/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1250 ALU_1b_0/comparator_0/AND_3/a_78_8# ALU_1b_0/AND_8/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 ALU_1b_0/comparator_0/NOR_2/A ALU_1b_0/comparator_0/AND_3/a_78_51# vdd ALU_1b_0/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1252 ALU_1b_0/comparator_0/AND_5/a_78_51# ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1253 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1254 vdd ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_5/a_78_51# ALU_1b_0/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1255 ALU_1b_0/comparator_0/AND_5/a_78_51# ALU_1b_0/AND_7/out vdd ALU_1b_0/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 ALU_1b_0/comparator_0/AND_5/a_78_8# ALU_1b_0/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_5/a_78_51# vdd ALU_1b_0/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1258 ALU_1b_0/comparator_0/AND_4/a_78_51# ALU_1b_0/AND_8/out ALU_1b_0/comparator_0/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1259 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1260 vdd ALU_1b_0/AND_8/out ALU_1b_0/comparator_0/AND_4/a_78_51# ALU_1b_0/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1261 ALU_1b_0/comparator_0/AND_4/a_78_51# ALU_1b_0/AND_7/out vdd ALU_1b_0/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1262 ALU_1b_0/comparator_0/AND_4/a_78_8# ALU_1b_0/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_4/a_78_51# vdd ALU_1b_0/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1264 gnd ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1265 ALU_1b_0/comparator_0/NOR_0/out ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/NOR_0/a_n14_7# ALU_1b_0/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1266 ALU_1b_0/comparator_0/NOR_0/a_n14_7# ALU_1b_0/comparator_0/NOR_0/A vdd ALU_1b_0/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 ALU_1b_0/comparator_0/NOR_0/out ALU_1b_0/comparator_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 gnd ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/comparator_0/NOR_1/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1269 ALU_1b_0/comparator_0/NOR_1/out ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/comparator_0/NOR_1/a_n14_7# ALU_1b_0/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1270 ALU_1b_0/comparator_0/NOR_1/a_n14_7# ALU_1b_0/comparator_0/NOR_1/A vdd ALU_1b_0/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 ALU_1b_0/comparator_0/NOR_1/out ALU_1b_0/comparator_0/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1272 vdd ALU_1b_0/comparator_0/NOR_1/out ALU_1b_0/AND_10/B ALU_1b_0/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1273 gnd ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_5/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1274 gnd ALU_1b_0/comparator_0/NOR_0/out ALU_1b_0/comparator_0/NOR_1/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1275 vdd ALU_1b_0/comparator_0/NOR_0/out ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1276 gnd ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/AND_11/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1277 vdd ALU_1b_0/comparator_0/NOR_3/out ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=9 ps=5
M1278 gnd ALU_1b_0/comparator_0/NOR_3/out ALU_1b_0/comparator_0/NOR_2/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1279 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1280 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/AND_7/out vdd ALU_1b_0/comparator_0/w_n39_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1281 gnd ALU_1b_0/comparator_0/NOR_1/out ALU_1b_0/AND_10/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1282 vdd ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/AND_11/B ALU_1b_0/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1283 vdd ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/w_n74_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=1 ps=1
M1284 ALU_1b_0/AND_19/A ALU_1b_0/NOT_1/in vdd ALU_1b_0/NOT_1/w_n36_43# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1285 ALU_1b_0/AND_19/A ALU_1b_0/NOT_1/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1286 ALU_1b_0/AND_3/A A0 vdd ALU_1b_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1287 ALU_1b_0/AND_3/A A0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1288 ALU_1b_0/NOR_2/A ALU_1b_0/NOT_2/in vdd ALU_1b_0/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1289 ALU_1b_0/NOR_2/A ALU_1b_0/NOT_2/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1290 ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/decoder_0/AND_1/B ALU_1b_0/decoder_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1291 ALU_1b_0/AND_2/B ALU_1b_0/decoder_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1292 vdd ALU_1b_0/decoder_0/AND_1/B ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1293 ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/decoder_0/AND_2/B vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 ALU_1b_0/decoder_0/AND_0/a_78_8# ALU_1b_0/decoder_0/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 ALU_1b_0/AND_2/B ALU_1b_0/decoder_0/AND_0/a_78_51# vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1296 ALU_1b_0/decoder_0/AND_1/a_78_51# ALU_1b_0/decoder_0/AND_1/B ALU_1b_0/decoder_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1297 ALU_1b_0/AND_9/A ALU_1b_0/decoder_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1298 vdd ALU_1b_0/decoder_0/AND_1/B ALU_1b_0/decoder_0/AND_1/a_78_51# ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1299 ALU_1b_0/decoder_0/AND_1/a_78_51# S1 vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 ALU_1b_0/decoder_0/AND_1/a_78_8# S1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1301 ALU_1b_0/AND_9/A ALU_1b_0/decoder_0/AND_1/a_78_51# vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1302 ALU_1b_0/decoder_0/AND_2/a_78_51# ALU_1b_0/decoder_0/AND_2/B ALU_1b_0/decoder_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1303 ALU_1b_0/AND_5/B ALU_1b_0/decoder_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1304 vdd ALU_1b_0/decoder_0/AND_2/B ALU_1b_0/decoder_0/AND_2/a_78_51# ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1305 ALU_1b_0/decoder_0/AND_2/a_78_51# S0 vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1306 ALU_1b_0/decoder_0/AND_2/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1307 ALU_1b_0/AND_5/B ALU_1b_0/decoder_0/AND_2/a_78_51# vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1308 ALU_1b_0/decoder_0/AND_3/a_78_51# S1 ALU_1b_0/decoder_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1309 ALU_1b_0/AND_15/A ALU_1b_0/decoder_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1310 vdd S1 ALU_1b_0/decoder_0/AND_3/a_78_51# ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1311 ALU_1b_0/decoder_0/AND_3/a_78_51# S0 vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 ALU_1b_0/decoder_0/AND_3/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1313 ALU_1b_0/AND_15/A ALU_1b_0/decoder_0/AND_3/a_78_51# vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1314 ALU_1b_0/decoder_0/AND_2/B S1 vdd ALU_1b_0/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1315 ALU_1b_0/decoder_0/AND_2/B S1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1316 ALU_1b_0/decoder_0/AND_1/B S0 vdd ALU_1b_0/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1317 ALU_1b_0/decoder_0/AND_1/B S0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1318 ALU_1b_0/NOR_2/B ALU_1b_0/NOT_3/in vdd ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1319 ALU_1b_0/NOR_2/B ALU_1b_0/NOT_3/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1320 gnd ALU_1b_0/NOR_0/B ALU_1b_0/NOT_2/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1321 ALU_1b_0/NOT_2/in ALU_1b_0/NOR_0/B ALU_1b_0/NOR_0/a_n14_7# ALU_1b_0/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1322 ALU_1b_0/NOR_0/a_n14_7# ALU_1b_0/NOR_0/A vdd ALU_1b_0/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 ALU_1b_0/NOT_2/in ALU_1b_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1324 F0 ALU_1b_0/NOT_4/in vdd ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1325 F0 ALU_1b_0/NOT_4/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1326 gnd ALU_1b_0/NOR_1/B ALU_1b_0/NOT_3/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1327 ALU_1b_0/NOT_3/in ALU_1b_0/NOR_1/B ALU_1b_0/NOR_1/a_n14_7# ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1328 ALU_1b_0/NOR_1/a_n14_7# ALU_1b_0/NOR_1/A vdd ALU_1b_0/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 ALU_1b_0/NOT_3/in ALU_1b_0/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1330 gnd ALU_1b_1/NOR_2/B ALU_1b_1/NOT_4/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1331 ALU_1b_1/NOT_4/in ALU_1b_1/NOR_2/B ALU_1b_1/NOR_2/a_n14_7# ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1332 ALU_1b_1/NOR_2/a_n14_7# ALU_1b_1/NOR_2/A vdd ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1333 ALU_1b_1/NOT_4/in ALU_1b_1/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 ALU_1b_1/NOR_4/B ALU_1b_1/NOT_5/in vdd ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1335 ALU_1b_1/NOR_4/B ALU_1b_1/NOT_5/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1336 Cout ALU_1b_1/NOT_6/in vdd ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1337 Cout ALU_1b_1/NOT_6/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1338 gnd ALU_1b_1/NOR_3/B ALU_1b_1/NOT_5/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1339 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_3/B ALU_1b_1/NOR_3/a_n14_7# ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1340 ALU_1b_1/NOR_3/a_n14_7# ALU_1b_1/NOR_3/A vdd ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1341 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1342 gnd ALU_1b_1/NOR_4/B ALU_1b_1/NOT_6/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1343 ALU_1b_1/NOT_6/in ALU_1b_1/NOR_4/B ALU_1b_1/NOR_4/a_n14_7# ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1344 ALU_1b_1/NOR_4/a_n14_7# ALU_1b_1/NOR_4/A vdd ALU_1b_1/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 ALU_1b_1/NOT_6/in ALU_1b_1/NOR_4/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1346 ALU_1b_1/AND_0/a_78_51# A3 ALU_1b_1/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1347 ALU_1b_1/AND_0/out ALU_1b_1/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1348 vdd A3 ALU_1b_1/AND_0/a_78_51# ALU_1b_1/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1349 ALU_1b_1/AND_0/a_78_51# ALU_1b_1/AND_2/B vdd ALU_1b_1/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1350 ALU_1b_1/AND_0/a_78_8# ALU_1b_1/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 ALU_1b_1/AND_0/out ALU_1b_1/AND_0/a_78_51# vdd ALU_1b_1/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1352 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1353 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out ALU_1b_1/full_adder_0/half_adder_1/A vdd ALU_1b_1/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1354 vdd ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out ALU_1b_1/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1355 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/a_n7_n34# ALU_1b_1/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1356 ALU_1b_1/AND_16/A ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1357 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_0/half_adder_1/A vdd ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1358 ALU_1b_1/AND_16/A ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1359 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_1/AND_1/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1360 gnd ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1361 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1362 vdd ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1363 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/AND_16/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_16/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 gnd ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1366 vdd ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1367 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1368 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out vdd ALU_1b_1/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1369 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1370 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1371 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out ALU_1b_1/AND_0/out vdd ALU_1b_1/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1372 vdd ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out ALU_1b_1/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1373 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_1/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1374 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1375 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_1/AND_0/out vdd ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1376 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1377 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# ALU_1b_1/AND_2/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1378 gnd ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1379 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 vdd ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1381 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_1/full_adder_0/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 gnd ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1384 vdd ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1385 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_1/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1386 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out vdd ALU_1b_1/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1387 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1388 gnd ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1389 ALU_1b_1/full_adder_0/NOR_0/out ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/NOR_0/a_n14_7# ALU_1b_1/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1390 ALU_1b_1/full_adder_0/NOR_0/a_n14_7# ALU_1b_1/full_adder_0/NOR_0/A vdd ALU_1b_1/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 ALU_1b_1/full_adder_0/NOR_0/out ALU_1b_1/full_adder_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1392 ALU_1b_1/AND_17/A ALU_1b_1/full_adder_0/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1393 ALU_1b_1/AND_17/A ALU_1b_1/full_adder_0/NOR_0/out vdd ALU_1b_1/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1394 ALU_1b_1/AND_1/a_78_51# ALU_1b_1/AND_2/B ALU_1b_1/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1395 ALU_1b_1/AND_1/out ALU_1b_1/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1396 vdd ALU_1b_1/AND_2/B ALU_1b_1/AND_1/a_78_51# ALU_1b_1/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1397 ALU_1b_1/AND_1/a_78_51# ALU_1b_1/C0 vdd ALU_1b_1/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1398 ALU_1b_1/AND_1/a_78_8# ALU_1b_1/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1399 ALU_1b_1/AND_1/out ALU_1b_1/AND_1/a_78_51# vdd ALU_1b_1/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1400 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1401 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/half_adder_1/A vdd ALU_1b_1/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1402 vdd ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/a_n7_n34# ALU_1b_1/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1404 ALU_1b_1/NOT_1/in ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1405 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_1/half_adder_1/A vdd ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1406 ALU_1b_1/NOT_1/in ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1407 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_1/AND_5/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1408 gnd ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1409 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 vdd ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1411 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_1/NOT_1/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/NOT_1/in ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1413 gnd ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1414 vdd ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1415 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1416 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out vdd ALU_1b_1/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1417 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1418 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1419 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/AND_3/out vdd ALU_1b_1/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1420 vdd ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1421 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_1/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1422 ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/AND_3/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1423 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_1/AND_3/out vdd ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1424 ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1425 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_1/AND_4/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1426 gnd ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1427 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 vdd ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1429 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_1/full_adder_1/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_1/AND_3/out ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 gnd ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1432 vdd ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1433 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_1/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1434 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out vdd ALU_1b_1/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1435 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1436 gnd ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1437 ALU_1b_1/full_adder_1/NOR_0/out ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/NOR_0/a_n14_7# ALU_1b_1/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1438 ALU_1b_1/full_adder_1/NOR_0/a_n14_7# ALU_1b_1/full_adder_1/NOR_0/A vdd ALU_1b_1/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1439 ALU_1b_1/full_adder_1/NOR_0/out ALU_1b_1/full_adder_1/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1440 ALU_1b_1/AND_18/A ALU_1b_1/full_adder_1/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1441 ALU_1b_1/AND_18/A ALU_1b_1/full_adder_1/NOR_0/out vdd ALU_1b_1/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1442 ALU_1b_1/AND_2/a_78_51# ALU_1b_1/AND_2/B ALU_1b_1/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1443 ALU_1b_1/AND_2/out ALU_1b_1/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1444 vdd ALU_1b_1/AND_2/B ALU_1b_1/AND_2/a_78_51# ALU_1b_1/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1445 ALU_1b_1/AND_2/a_78_51# B3 vdd ALU_1b_1/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 ALU_1b_1/AND_2/a_78_8# B3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 ALU_1b_1/AND_2/out ALU_1b_1/AND_2/a_78_51# vdd ALU_1b_1/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1448 ALU_1b_1/AND_3/a_78_51# ALU_1b_1/AND_5/B ALU_1b_1/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1449 ALU_1b_1/AND_3/out ALU_1b_1/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1450 vdd ALU_1b_1/AND_5/B ALU_1b_1/AND_3/a_78_51# ALU_1b_1/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1451 ALU_1b_1/AND_3/a_78_51# ALU_1b_1/AND_3/A vdd ALU_1b_1/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 ALU_1b_1/AND_3/a_78_8# ALU_1b_1/AND_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 ALU_1b_1/AND_3/out ALU_1b_1/AND_3/a_78_51# vdd ALU_1b_1/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1454 ALU_1b_1/AND_5/a_78_51# ALU_1b_1/AND_5/B ALU_1b_1/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1455 ALU_1b_1/AND_5/out ALU_1b_1/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1456 vdd ALU_1b_1/AND_5/B ALU_1b_1/AND_5/a_78_51# ALU_1b_1/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1457 ALU_1b_1/AND_5/a_78_51# ALU_1b_1/C0 vdd ALU_1b_1/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1458 ALU_1b_1/AND_5/a_78_8# ALU_1b_1/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1459 ALU_1b_1/AND_5/out ALU_1b_1/AND_5/a_78_51# vdd ALU_1b_1/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1460 ALU_1b_1/AND_4/a_78_51# ALU_1b_1/AND_5/B ALU_1b_1/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1461 ALU_1b_1/AND_4/out ALU_1b_1/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1462 vdd ALU_1b_1/AND_5/B ALU_1b_1/AND_4/a_78_51# ALU_1b_1/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1463 ALU_1b_1/AND_4/a_78_51# B3 vdd ALU_1b_1/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1464 ALU_1b_1/AND_4/a_78_8# B3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 ALU_1b_1/AND_4/out ALU_1b_1/AND_4/a_78_51# vdd ALU_1b_1/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1466 ALU_1b_1/AND_10/a_78_51# ALU_1b_1/AND_10/B ALU_1b_1/AND_10/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1467 ALU_1b_1/NOR_1/A ALU_1b_1/AND_10/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1468 vdd ALU_1b_1/AND_10/B ALU_1b_1/AND_10/a_78_51# ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1469 ALU_1b_1/AND_10/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1470 ALU_1b_1/AND_10/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1471 ALU_1b_1/NOR_1/A ALU_1b_1/AND_10/a_78_51# vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1472 ALU_1b_1/AND_11/a_78_51# ALU_1b_1/AND_11/B ALU_1b_1/AND_11/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1473 ALU_1b_1/NOR_4/A ALU_1b_1/AND_11/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1474 vdd ALU_1b_1/AND_11/B ALU_1b_1/AND_11/a_78_51# ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1475 ALU_1b_1/AND_11/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 ALU_1b_1/AND_11/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1477 ALU_1b_1/NOR_4/A ALU_1b_1/AND_11/a_78_51# vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1478 ALU_1b_1/AND_6/a_78_51# A3 ALU_1b_1/AND_6/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1479 ALU_1b_1/AND_6/out ALU_1b_1/AND_6/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1480 vdd A3 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1481 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 ALU_1b_1/AND_6/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1483 ALU_1b_1/AND_6/out ALU_1b_1/AND_6/a_78_51# vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1484 ALU_1b_1/AND_7/a_78_51# B3 ALU_1b_1/AND_7/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1485 ALU_1b_1/AND_7/out ALU_1b_1/AND_7/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1486 vdd B3 ALU_1b_1/AND_7/a_78_51# ALU_1b_1/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1487 ALU_1b_1/AND_7/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 ALU_1b_1/AND_7/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 ALU_1b_1/AND_7/out ALU_1b_1/AND_7/a_78_51# vdd ALU_1b_1/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1490 ALU_1b_1/AND_12/a_78_51# A3 ALU_1b_1/AND_12/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1491 ALU_1b_1/AND_14/B ALU_1b_1/AND_12/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1492 vdd A3 ALU_1b_1/AND_12/a_78_51# ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1493 ALU_1b_1/AND_12/a_78_51# ALU_1b_1/AND_15/A vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 ALU_1b_1/AND_12/a_78_8# ALU_1b_1/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1495 ALU_1b_1/AND_14/B ALU_1b_1/AND_12/a_78_51# vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1496 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/C0 ALU_1b_1/AND_8/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1497 ALU_1b_1/AND_8/out ALU_1b_1/AND_8/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1498 vdd ALU_1b_1/C0 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1499 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1500 ALU_1b_1/AND_8/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1501 ALU_1b_1/AND_8/out ALU_1b_1/AND_8/a_78_51# vdd ALU_1b_1/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1502 ALU_1b_1/AND_13/a_78_51# B3 ALU_1b_1/AND_13/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1503 ALU_1b_1/AND_14/A ALU_1b_1/AND_13/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1504 vdd B3 ALU_1b_1/AND_13/a_78_51# ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1505 ALU_1b_1/AND_13/a_78_51# ALU_1b_1/AND_15/A vdd ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1506 ALU_1b_1/AND_13/a_78_8# ALU_1b_1/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1507 ALU_1b_1/AND_14/A ALU_1b_1/AND_13/a_78_51# vdd ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1508 ALU_1b_1/AND_9/a_78_51# F2 ALU_1b_1/AND_9/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1509 ALU_1b_1/AND_9/out ALU_1b_1/AND_9/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1510 vdd F2 ALU_1b_1/AND_9/a_78_51# ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1511 ALU_1b_1/AND_9/a_78_51# ALU_1b_1/AND_9/A vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1512 ALU_1b_1/AND_9/a_78_8# ALU_1b_1/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1513 ALU_1b_1/AND_9/out ALU_1b_1/AND_9/a_78_51# vdd ALU_1b_1/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1514 ALU_1b_1/AND_14/a_78_51# ALU_1b_1/AND_14/B ALU_1b_1/AND_14/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1515 ALU_1b_1/AND_15/B ALU_1b_1/AND_14/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1516 vdd ALU_1b_1/AND_14/B ALU_1b_1/AND_14/a_78_51# ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1517 ALU_1b_1/AND_14/a_78_51# ALU_1b_1/AND_14/A vdd ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 ALU_1b_1/AND_14/a_78_8# ALU_1b_1/AND_14/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1519 ALU_1b_1/AND_15/B ALU_1b_1/AND_14/a_78_51# vdd ALU_1b_1/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1520 ALU_1b_1/AND_15/a_78_51# ALU_1b_1/AND_15/B ALU_1b_1/AND_15/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1521 ALU_1b_1/NOR_1/B ALU_1b_1/AND_15/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1522 vdd ALU_1b_1/AND_15/B ALU_1b_1/AND_15/a_78_51# ALU_1b_1/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1523 ALU_1b_1/AND_15/a_78_51# ALU_1b_1/AND_15/A vdd ALU_1b_1/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 ALU_1b_1/AND_15/a_78_8# ALU_1b_1/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 ALU_1b_1/NOR_1/B ALU_1b_1/AND_15/a_78_51# vdd ALU_1b_1/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1526 ALU_1b_1/AND_16/a_78_51# ALU_1b_1/AND_2/B ALU_1b_1/AND_16/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1527 ALU_1b_1/NOR_0/B ALU_1b_1/AND_16/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1528 vdd ALU_1b_1/AND_2/B ALU_1b_1/AND_16/a_78_51# ALU_1b_1/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1529 ALU_1b_1/AND_16/a_78_51# ALU_1b_1/AND_16/A vdd ALU_1b_1/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1530 ALU_1b_1/AND_16/a_78_8# ALU_1b_1/AND_16/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 ALU_1b_1/NOR_0/B ALU_1b_1/AND_16/a_78_51# vdd ALU_1b_1/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1532 ALU_1b_1/AND_17/a_78_51# ALU_1b_1/AND_2/B ALU_1b_1/AND_17/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1533 ALU_1b_1/NOR_3/B ALU_1b_1/AND_17/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1534 vdd ALU_1b_1/AND_2/B ALU_1b_1/AND_17/a_78_51# ALU_1b_1/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1535 ALU_1b_1/AND_17/a_78_51# ALU_1b_1/AND_17/A vdd ALU_1b_1/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 ALU_1b_1/AND_17/a_78_8# ALU_1b_1/AND_17/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 ALU_1b_1/NOR_3/B ALU_1b_1/AND_17/a_78_51# vdd ALU_1b_1/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1538 ALU_1b_1/AND_19/a_78_51# ALU_1b_1/AND_5/B ALU_1b_1/AND_19/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1539 ALU_1b_1/NOR_0/A ALU_1b_1/AND_19/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1540 vdd ALU_1b_1/AND_5/B ALU_1b_1/AND_19/a_78_51# ALU_1b_1/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1541 ALU_1b_1/AND_19/a_78_51# ALU_1b_1/AND_19/A vdd ALU_1b_1/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1542 ALU_1b_1/AND_19/a_78_8# ALU_1b_1/AND_19/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1543 ALU_1b_1/NOR_0/A ALU_1b_1/AND_19/a_78_51# vdd ALU_1b_1/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1544 ALU_1b_1/AND_18/a_78_51# ALU_1b_1/AND_5/B ALU_1b_1/AND_18/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1545 ALU_1b_1/NOR_3/A ALU_1b_1/AND_18/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1546 vdd ALU_1b_1/AND_5/B ALU_1b_1/AND_18/a_78_51# ALU_1b_1/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1547 ALU_1b_1/AND_18/a_78_51# ALU_1b_1/AND_18/A vdd ALU_1b_1/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1548 ALU_1b_1/AND_18/a_78_8# ALU_1b_1/AND_18/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 ALU_1b_1/NOR_3/A ALU_1b_1/AND_18/a_78_51# vdd ALU_1b_1/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1550 gnd ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_2/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1551 ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_2/a_n14_7# ALU_1b_1/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1552 ALU_1b_1/comparator_0/NOR_2/a_n14_7# ALU_1b_1/comparator_0/NOR_2/A vdd ALU_1b_1/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1553 ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/comparator_0/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1554 gnd ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/NOR_3/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1555 ALU_1b_1/comparator_0/NOR_3/out ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/NOR_3/a_n14_7# ALU_1b_1/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1556 ALU_1b_1/comparator_0/NOR_3/a_n14_7# ALU_1b_1/comparator_0/NOR_3/A vdd ALU_1b_1/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 ALU_1b_1/comparator_0/NOR_3/out ALU_1b_1/comparator_0/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 ALU_1b_1/comparator_0/AND_0/a_78_51# ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1559 ALU_1b_1/comparator_0/NOR_0/A ALU_1b_1/comparator_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1560 vdd ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_0/a_78_51# ALU_1b_1/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1561 ALU_1b_1/comparator_0/AND_0/a_78_51# ALU_1b_1/AND_6/out vdd ALU_1b_1/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1562 ALU_1b_1/comparator_0/AND_0/a_78_8# ALU_1b_1/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1563 ALU_1b_1/comparator_0/NOR_0/A ALU_1b_1/comparator_0/AND_0/a_78_51# vdd ALU_1b_1/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1564 ALU_1b_1/comparator_0/AND_1/a_78_51# ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1565 ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1566 vdd ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/AND_1/a_78_51# ALU_1b_1/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1567 ALU_1b_1/comparator_0/AND_1/a_78_51# ALU_1b_1/AND_6/out vdd ALU_1b_1/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1568 ALU_1b_1/comparator_0/AND_1/a_78_8# ALU_1b_1/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1569 ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/AND_1/a_78_51# vdd ALU_1b_1/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1570 ALU_1b_1/comparator_0/AND_2/a_78_51# ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1571 ALU_1b_1/comparator_0/NOR_1/A ALU_1b_1/comparator_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1572 vdd ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_2/a_78_51# ALU_1b_1/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1573 ALU_1b_1/comparator_0/AND_2/a_78_51# ALU_1b_1/AND_9/out vdd ALU_1b_1/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1574 ALU_1b_1/comparator_0/AND_2/a_78_8# ALU_1b_1/AND_9/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1575 ALU_1b_1/comparator_0/NOR_1/A ALU_1b_1/comparator_0/AND_2/a_78_51# vdd ALU_1b_1/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1576 ALU_1b_1/comparator_0/AND_3/a_78_51# ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1577 ALU_1b_1/comparator_0/NOR_2/A ALU_1b_1/comparator_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1578 vdd ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_3/a_78_51# ALU_1b_1/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1579 ALU_1b_1/comparator_0/AND_3/a_78_51# ALU_1b_1/AND_8/out vdd ALU_1b_1/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1580 ALU_1b_1/comparator_0/AND_3/a_78_8# ALU_1b_1/AND_8/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1581 ALU_1b_1/comparator_0/NOR_2/A ALU_1b_1/comparator_0/AND_3/a_78_51# vdd ALU_1b_1/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1582 ALU_1b_1/comparator_0/AND_5/a_78_51# ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1583 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1584 vdd ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_5/a_78_51# ALU_1b_1/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1585 ALU_1b_1/comparator_0/AND_5/a_78_51# ALU_1b_1/AND_7/out vdd ALU_1b_1/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1586 ALU_1b_1/comparator_0/AND_5/a_78_8# ALU_1b_1/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1587 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_5/a_78_51# vdd ALU_1b_1/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1588 ALU_1b_1/comparator_0/AND_4/a_78_51# ALU_1b_1/AND_8/out ALU_1b_1/comparator_0/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1589 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1590 vdd ALU_1b_1/AND_8/out ALU_1b_1/comparator_0/AND_4/a_78_51# ALU_1b_1/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1591 ALU_1b_1/comparator_0/AND_4/a_78_51# ALU_1b_1/AND_7/out vdd ALU_1b_1/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 ALU_1b_1/comparator_0/AND_4/a_78_8# ALU_1b_1/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_4/a_78_51# vdd ALU_1b_1/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1594 gnd ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1595 ALU_1b_1/comparator_0/NOR_0/out ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/NOR_0/a_n14_7# ALU_1b_1/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1596 ALU_1b_1/comparator_0/NOR_0/a_n14_7# ALU_1b_1/comparator_0/NOR_0/A vdd ALU_1b_1/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 ALU_1b_1/comparator_0/NOR_0/out ALU_1b_1/comparator_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1598 gnd ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/comparator_0/NOR_1/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1599 ALU_1b_1/comparator_0/NOR_1/out ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/comparator_0/NOR_1/a_n14_7# ALU_1b_1/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1600 ALU_1b_1/comparator_0/NOR_1/a_n14_7# ALU_1b_1/comparator_0/NOR_1/A vdd ALU_1b_1/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1601 ALU_1b_1/comparator_0/NOR_1/out ALU_1b_1/comparator_0/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1602 vdd ALU_1b_1/comparator_0/NOR_1/out ALU_1b_1/AND_10/B ALU_1b_1/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1603 gnd ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_5/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1604 gnd ALU_1b_1/comparator_0/NOR_0/out ALU_1b_1/comparator_0/NOR_1/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1605 vdd ALU_1b_1/comparator_0/NOR_0/out ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1606 gnd ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/AND_11/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1607 vdd ALU_1b_1/comparator_0/NOR_3/out ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=9 ps=5
M1608 gnd ALU_1b_1/comparator_0/NOR_3/out ALU_1b_1/comparator_0/NOR_2/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1609 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1610 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/AND_7/out vdd ALU_1b_1/comparator_0/w_n39_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1611 gnd ALU_1b_1/comparator_0/NOR_1/out ALU_1b_1/AND_10/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1612 vdd ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/AND_11/B ALU_1b_1/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1613 vdd ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/w_n74_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=1 ps=1
M1614 ALU_1b_1/AND_19/A ALU_1b_1/NOT_1/in vdd ALU_1b_1/NOT_1/w_n36_43# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1615 ALU_1b_1/AND_19/A ALU_1b_1/NOT_1/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1616 ALU_1b_1/AND_3/A A3 vdd ALU_1b_1/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1617 ALU_1b_1/AND_3/A A3 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1618 ALU_1b_1/NOR_2/A ALU_1b_1/NOT_2/in vdd ALU_1b_1/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1619 ALU_1b_1/NOR_2/A ALU_1b_1/NOT_2/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1620 ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/decoder_0/AND_1/B ALU_1b_1/decoder_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1621 ALU_1b_1/AND_2/B ALU_1b_1/decoder_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1622 vdd ALU_1b_1/decoder_0/AND_1/B ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1623 ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/decoder_0/AND_2/B vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1624 ALU_1b_1/decoder_0/AND_0/a_78_8# ALU_1b_1/decoder_0/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 ALU_1b_1/AND_2/B ALU_1b_1/decoder_0/AND_0/a_78_51# vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1626 ALU_1b_1/decoder_0/AND_1/a_78_51# ALU_1b_1/decoder_0/AND_1/B ALU_1b_1/decoder_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1627 ALU_1b_1/AND_9/A ALU_1b_1/decoder_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1628 vdd ALU_1b_1/decoder_0/AND_1/B ALU_1b_1/decoder_0/AND_1/a_78_51# ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1629 ALU_1b_1/decoder_0/AND_1/a_78_51# S1 vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1630 ALU_1b_1/decoder_0/AND_1/a_78_8# S1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1631 ALU_1b_1/AND_9/A ALU_1b_1/decoder_0/AND_1/a_78_51# vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1632 ALU_1b_1/decoder_0/AND_2/a_78_51# ALU_1b_1/decoder_0/AND_2/B ALU_1b_1/decoder_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1633 ALU_1b_1/AND_5/B ALU_1b_1/decoder_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1634 vdd ALU_1b_1/decoder_0/AND_2/B ALU_1b_1/decoder_0/AND_2/a_78_51# ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1635 ALU_1b_1/decoder_0/AND_2/a_78_51# S0 vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1636 ALU_1b_1/decoder_0/AND_2/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 ALU_1b_1/AND_5/B ALU_1b_1/decoder_0/AND_2/a_78_51# vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1638 ALU_1b_1/decoder_0/AND_3/a_78_51# S1 ALU_1b_1/decoder_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1639 ALU_1b_1/AND_15/A ALU_1b_1/decoder_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1640 vdd S1 ALU_1b_1/decoder_0/AND_3/a_78_51# ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1641 ALU_1b_1/decoder_0/AND_3/a_78_51# S0 vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1642 ALU_1b_1/decoder_0/AND_3/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1643 ALU_1b_1/AND_15/A ALU_1b_1/decoder_0/AND_3/a_78_51# vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1644 ALU_1b_1/decoder_0/AND_2/B S1 vdd ALU_1b_1/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1645 ALU_1b_1/decoder_0/AND_2/B S1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1646 ALU_1b_1/decoder_0/AND_1/B S0 vdd ALU_1b_1/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1647 ALU_1b_1/decoder_0/AND_1/B S0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1648 ALU_1b_1/NOR_2/B ALU_1b_1/NOT_3/in vdd ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1649 ALU_1b_1/NOR_2/B ALU_1b_1/NOT_3/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1650 gnd ALU_1b_1/NOR_0/B ALU_1b_1/NOT_2/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1651 ALU_1b_1/NOT_2/in ALU_1b_1/NOR_0/B ALU_1b_1/NOR_0/a_n14_7# ALU_1b_1/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1652 ALU_1b_1/NOR_0/a_n14_7# ALU_1b_1/NOR_0/A vdd ALU_1b_1/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1653 ALU_1b_1/NOT_2/in ALU_1b_1/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1654 F3 ALU_1b_1/NOT_4/in vdd ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1655 F3 ALU_1b_1/NOT_4/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1656 gnd ALU_1b_1/NOR_1/B ALU_1b_1/NOT_3/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1657 ALU_1b_1/NOT_3/in ALU_1b_1/NOR_1/B ALU_1b_1/NOR_1/a_n14_7# ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1658 ALU_1b_1/NOR_1/a_n14_7# ALU_1b_1/NOR_1/A vdd ALU_1b_1/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1659 ALU_1b_1/NOT_3/in ALU_1b_1/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1660 gnd ALU_1b_2/NOR_2/B ALU_1b_2/NOT_4/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1661 ALU_1b_2/NOT_4/in ALU_1b_2/NOR_2/B ALU_1b_2/NOR_2/a_n14_7# ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1662 ALU_1b_2/NOR_2/a_n14_7# ALU_1b_2/NOR_2/A vdd ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1663 ALU_1b_2/NOT_4/in ALU_1b_2/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 ALU_1b_2/NOR_4/B ALU_1b_2/NOT_5/in vdd ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1665 ALU_1b_2/NOR_4/B ALU_1b_2/NOT_5/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1666 ALU_1b_3/C0 ALU_1b_2/NOT_6/in vdd ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1667 ALU_1b_3/C0 ALU_1b_2/NOT_6/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1668 gnd ALU_1b_2/NOR_3/B ALU_1b_2/NOT_5/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1669 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_3/B ALU_1b_2/NOR_3/a_n14_7# ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1670 ALU_1b_2/NOR_3/a_n14_7# ALU_1b_2/NOR_3/A vdd ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1671 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1672 gnd ALU_1b_2/NOR_4/B ALU_1b_2/NOT_6/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1673 ALU_1b_2/NOT_6/in ALU_1b_2/NOR_4/B ALU_1b_2/NOR_4/a_n14_7# ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1674 ALU_1b_2/NOR_4/a_n14_7# ALU_1b_2/NOR_4/A vdd ALU_1b_2/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1675 ALU_1b_2/NOT_6/in ALU_1b_2/NOR_4/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1676 ALU_1b_2/AND_0/a_78_51# A1 ALU_1b_2/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1677 ALU_1b_2/AND_0/out ALU_1b_2/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1678 vdd A1 ALU_1b_2/AND_0/a_78_51# ALU_1b_2/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1679 ALU_1b_2/AND_0/a_78_51# ALU_1b_2/AND_2/B vdd ALU_1b_2/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 ALU_1b_2/AND_0/a_78_8# ALU_1b_2/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 ALU_1b_2/AND_0/out ALU_1b_2/AND_0/a_78_51# vdd ALU_1b_2/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1682 ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1683 ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out ALU_1b_2/full_adder_0/half_adder_1/A vdd ALU_1b_2/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1684 vdd ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out ALU_1b_2/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 ALU_1b_2/full_adder_0/half_adder_1/NAND_0/a_n7_n34# ALU_1b_2/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1686 ALU_1b_2/AND_16/A ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1687 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_0/half_adder_1/A vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1688 ALU_1b_2/AND_16/A ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1689 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_2/AND_1/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1690 gnd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1691 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1692 vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1693 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/AND_16/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1694 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_16/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1695 gnd ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1696 vdd ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1697 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1698 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out vdd ALU_1b_2/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1699 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1700 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1701 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out ALU_1b_2/AND_0/out vdd ALU_1b_2/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1702 vdd ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out ALU_1b_2/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1703 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_2/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1704 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1705 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_2/AND_0/out vdd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1706 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1707 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# ALU_1b_2/AND_2/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1708 gnd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1709 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1710 vdd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1711 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_2/full_adder_0/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1712 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1713 gnd ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1714 vdd ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1715 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_2/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1716 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out vdd ALU_1b_2/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1717 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1718 gnd ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1719 ALU_1b_2/full_adder_0/NOR_0/out ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/NOR_0/a_n14_7# ALU_1b_2/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1720 ALU_1b_2/full_adder_0/NOR_0/a_n14_7# ALU_1b_2/full_adder_0/NOR_0/A vdd ALU_1b_2/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1721 ALU_1b_2/full_adder_0/NOR_0/out ALU_1b_2/full_adder_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1722 ALU_1b_2/AND_17/A ALU_1b_2/full_adder_0/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1723 ALU_1b_2/AND_17/A ALU_1b_2/full_adder_0/NOR_0/out vdd ALU_1b_2/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1724 ALU_1b_2/AND_1/a_78_51# ALU_1b_2/AND_2/B ALU_1b_2/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1725 ALU_1b_2/AND_1/out ALU_1b_2/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1726 vdd ALU_1b_2/AND_2/B ALU_1b_2/AND_1/a_78_51# ALU_1b_2/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1727 ALU_1b_2/AND_1/a_78_51# ALU_1b_2/C0 vdd ALU_1b_2/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1728 ALU_1b_2/AND_1/a_78_8# ALU_1b_2/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 ALU_1b_2/AND_1/out ALU_1b_2/AND_1/a_78_51# vdd ALU_1b_2/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1730 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1731 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/full_adder_1/half_adder_1/A vdd ALU_1b_2/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1732 vdd ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/a_n7_n34# ALU_1b_2/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1734 ALU_1b_2/NOT_1/in ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1735 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_1/half_adder_1/A vdd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1736 ALU_1b_2/NOT_1/in ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1737 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_2/AND_5/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1738 gnd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1739 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1740 vdd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1741 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_2/NOT_1/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1742 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/NOT_1/in ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1743 gnd ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1744 vdd ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1745 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1746 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out vdd ALU_1b_2/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1747 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1748 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1749 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/AND_3/out vdd ALU_1b_2/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1750 vdd ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1751 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_2/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1752 ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/AND_3/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1753 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_2/AND_3/out vdd ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1754 ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1755 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_2/AND_4/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1756 gnd ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1757 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1758 vdd ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1759 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_2/full_adder_1/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1760 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_2/AND_3/out ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1761 gnd ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1762 vdd ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1763 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_2/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1764 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out vdd ALU_1b_2/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1765 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1766 gnd ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1767 ALU_1b_2/full_adder_1/NOR_0/out ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/NOR_0/a_n14_7# ALU_1b_2/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1768 ALU_1b_2/full_adder_1/NOR_0/a_n14_7# ALU_1b_2/full_adder_1/NOR_0/A vdd ALU_1b_2/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1769 ALU_1b_2/full_adder_1/NOR_0/out ALU_1b_2/full_adder_1/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1770 ALU_1b_2/AND_18/A ALU_1b_2/full_adder_1/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1771 ALU_1b_2/AND_18/A ALU_1b_2/full_adder_1/NOR_0/out vdd ALU_1b_2/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1772 ALU_1b_2/AND_2/a_78_51# ALU_1b_2/AND_2/B ALU_1b_2/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1773 ALU_1b_2/AND_2/out ALU_1b_2/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1774 vdd ALU_1b_2/AND_2/B ALU_1b_2/AND_2/a_78_51# ALU_1b_2/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1775 ALU_1b_2/AND_2/a_78_51# B1 vdd ALU_1b_2/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1776 ALU_1b_2/AND_2/a_78_8# B1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1777 ALU_1b_2/AND_2/out ALU_1b_2/AND_2/a_78_51# vdd ALU_1b_2/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1778 ALU_1b_2/AND_3/a_78_51# ALU_1b_2/AND_5/B ALU_1b_2/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1779 ALU_1b_2/AND_3/out ALU_1b_2/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1780 vdd ALU_1b_2/AND_5/B ALU_1b_2/AND_3/a_78_51# ALU_1b_2/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1781 ALU_1b_2/AND_3/a_78_51# ALU_1b_2/AND_3/A vdd ALU_1b_2/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1782 ALU_1b_2/AND_3/a_78_8# ALU_1b_2/AND_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1783 ALU_1b_2/AND_3/out ALU_1b_2/AND_3/a_78_51# vdd ALU_1b_2/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1784 ALU_1b_2/AND_5/a_78_51# ALU_1b_2/AND_5/B ALU_1b_2/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1785 ALU_1b_2/AND_5/out ALU_1b_2/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1786 vdd ALU_1b_2/AND_5/B ALU_1b_2/AND_5/a_78_51# ALU_1b_2/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1787 ALU_1b_2/AND_5/a_78_51# ALU_1b_2/C0 vdd ALU_1b_2/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1788 ALU_1b_2/AND_5/a_78_8# ALU_1b_2/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1789 ALU_1b_2/AND_5/out ALU_1b_2/AND_5/a_78_51# vdd ALU_1b_2/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1790 ALU_1b_2/AND_4/a_78_51# ALU_1b_2/AND_5/B ALU_1b_2/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1791 ALU_1b_2/AND_4/out ALU_1b_2/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1792 vdd ALU_1b_2/AND_5/B ALU_1b_2/AND_4/a_78_51# ALU_1b_2/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1793 ALU_1b_2/AND_4/a_78_51# B1 vdd ALU_1b_2/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1794 ALU_1b_2/AND_4/a_78_8# B1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1795 ALU_1b_2/AND_4/out ALU_1b_2/AND_4/a_78_51# vdd ALU_1b_2/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1796 ALU_1b_2/AND_10/a_78_51# ALU_1b_2/AND_10/B ALU_1b_2/AND_10/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1797 ALU_1b_2/NOR_1/A ALU_1b_2/AND_10/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1798 vdd ALU_1b_2/AND_10/B ALU_1b_2/AND_10/a_78_51# ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1799 ALU_1b_2/AND_10/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1800 ALU_1b_2/AND_10/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1801 ALU_1b_2/NOR_1/A ALU_1b_2/AND_10/a_78_51# vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1802 ALU_1b_2/AND_11/a_78_51# ALU_1b_2/AND_11/B ALU_1b_2/AND_11/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1803 ALU_1b_2/NOR_4/A ALU_1b_2/AND_11/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1804 vdd ALU_1b_2/AND_11/B ALU_1b_2/AND_11/a_78_51# ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1805 ALU_1b_2/AND_11/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1806 ALU_1b_2/AND_11/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1807 ALU_1b_2/NOR_4/A ALU_1b_2/AND_11/a_78_51# vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1808 ALU_1b_2/AND_6/a_78_51# A1 ALU_1b_2/AND_6/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1809 ALU_1b_2/AND_6/out ALU_1b_2/AND_6/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1810 vdd A1 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1811 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1812 ALU_1b_2/AND_6/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1813 ALU_1b_2/AND_6/out ALU_1b_2/AND_6/a_78_51# vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1814 ALU_1b_2/AND_7/a_78_51# B1 ALU_1b_2/AND_7/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1815 ALU_1b_2/AND_7/out ALU_1b_2/AND_7/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1816 vdd B1 ALU_1b_2/AND_7/a_78_51# ALU_1b_2/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1817 ALU_1b_2/AND_7/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1818 ALU_1b_2/AND_7/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1819 ALU_1b_2/AND_7/out ALU_1b_2/AND_7/a_78_51# vdd ALU_1b_2/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1820 ALU_1b_2/AND_12/a_78_51# A1 ALU_1b_2/AND_12/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1821 ALU_1b_2/AND_14/B ALU_1b_2/AND_12/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1822 vdd A1 ALU_1b_2/AND_12/a_78_51# ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1823 ALU_1b_2/AND_12/a_78_51# ALU_1b_2/AND_15/A vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1824 ALU_1b_2/AND_12/a_78_8# ALU_1b_2/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1825 ALU_1b_2/AND_14/B ALU_1b_2/AND_12/a_78_51# vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1826 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/C0 ALU_1b_2/AND_8/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1827 ALU_1b_2/AND_8/out ALU_1b_2/AND_8/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1828 vdd ALU_1b_2/C0 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1829 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1830 ALU_1b_2/AND_8/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1831 ALU_1b_2/AND_8/out ALU_1b_2/AND_8/a_78_51# vdd ALU_1b_2/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1832 ALU_1b_2/AND_13/a_78_51# B1 ALU_1b_2/AND_13/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1833 ALU_1b_2/AND_14/A ALU_1b_2/AND_13/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1834 vdd B1 ALU_1b_2/AND_13/a_78_51# ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1835 ALU_1b_2/AND_13/a_78_51# ALU_1b_2/AND_15/A vdd ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1836 ALU_1b_2/AND_13/a_78_8# ALU_1b_2/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1837 ALU_1b_2/AND_14/A ALU_1b_2/AND_13/a_78_51# vdd ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1838 ALU_1b_2/AND_9/a_78_51# F0 ALU_1b_2/AND_9/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1839 ALU_1b_2/AND_9/out ALU_1b_2/AND_9/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1840 vdd F0 ALU_1b_2/AND_9/a_78_51# ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1841 ALU_1b_2/AND_9/a_78_51# ALU_1b_2/AND_9/A vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1842 ALU_1b_2/AND_9/a_78_8# ALU_1b_2/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1843 ALU_1b_2/AND_9/out ALU_1b_2/AND_9/a_78_51# vdd ALU_1b_2/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1844 ALU_1b_2/AND_14/a_78_51# ALU_1b_2/AND_14/B ALU_1b_2/AND_14/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1845 ALU_1b_2/AND_15/B ALU_1b_2/AND_14/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1846 vdd ALU_1b_2/AND_14/B ALU_1b_2/AND_14/a_78_51# ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1847 ALU_1b_2/AND_14/a_78_51# ALU_1b_2/AND_14/A vdd ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1848 ALU_1b_2/AND_14/a_78_8# ALU_1b_2/AND_14/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1849 ALU_1b_2/AND_15/B ALU_1b_2/AND_14/a_78_51# vdd ALU_1b_2/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1850 ALU_1b_2/AND_15/a_78_51# ALU_1b_2/AND_15/B ALU_1b_2/AND_15/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1851 ALU_1b_2/NOR_1/B ALU_1b_2/AND_15/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1852 vdd ALU_1b_2/AND_15/B ALU_1b_2/AND_15/a_78_51# ALU_1b_2/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1853 ALU_1b_2/AND_15/a_78_51# ALU_1b_2/AND_15/A vdd ALU_1b_2/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1854 ALU_1b_2/AND_15/a_78_8# ALU_1b_2/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1855 ALU_1b_2/NOR_1/B ALU_1b_2/AND_15/a_78_51# vdd ALU_1b_2/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1856 ALU_1b_2/AND_16/a_78_51# ALU_1b_2/AND_2/B ALU_1b_2/AND_16/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1857 ALU_1b_2/NOR_0/B ALU_1b_2/AND_16/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1858 vdd ALU_1b_2/AND_2/B ALU_1b_2/AND_16/a_78_51# ALU_1b_2/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1859 ALU_1b_2/AND_16/a_78_51# ALU_1b_2/AND_16/A vdd ALU_1b_2/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1860 ALU_1b_2/AND_16/a_78_8# ALU_1b_2/AND_16/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1861 ALU_1b_2/NOR_0/B ALU_1b_2/AND_16/a_78_51# vdd ALU_1b_2/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1862 ALU_1b_2/AND_17/a_78_51# ALU_1b_2/AND_2/B ALU_1b_2/AND_17/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1863 ALU_1b_2/NOR_3/B ALU_1b_2/AND_17/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1864 vdd ALU_1b_2/AND_2/B ALU_1b_2/AND_17/a_78_51# ALU_1b_2/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1865 ALU_1b_2/AND_17/a_78_51# ALU_1b_2/AND_17/A vdd ALU_1b_2/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1866 ALU_1b_2/AND_17/a_78_8# ALU_1b_2/AND_17/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1867 ALU_1b_2/NOR_3/B ALU_1b_2/AND_17/a_78_51# vdd ALU_1b_2/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1868 ALU_1b_2/AND_19/a_78_51# ALU_1b_2/AND_5/B ALU_1b_2/AND_19/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1869 ALU_1b_2/NOR_0/A ALU_1b_2/AND_19/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1870 vdd ALU_1b_2/AND_5/B ALU_1b_2/AND_19/a_78_51# ALU_1b_2/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1871 ALU_1b_2/AND_19/a_78_51# ALU_1b_2/AND_19/A vdd ALU_1b_2/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 ALU_1b_2/AND_19/a_78_8# ALU_1b_2/AND_19/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1873 ALU_1b_2/NOR_0/A ALU_1b_2/AND_19/a_78_51# vdd ALU_1b_2/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1874 ALU_1b_2/AND_18/a_78_51# ALU_1b_2/AND_5/B ALU_1b_2/AND_18/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1875 ALU_1b_2/NOR_3/A ALU_1b_2/AND_18/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1876 vdd ALU_1b_2/AND_5/B ALU_1b_2/AND_18/a_78_51# ALU_1b_2/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1877 ALU_1b_2/AND_18/a_78_51# ALU_1b_2/AND_18/A vdd ALU_1b_2/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1878 ALU_1b_2/AND_18/a_78_8# ALU_1b_2/AND_18/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1879 ALU_1b_2/NOR_3/A ALU_1b_2/AND_18/a_78_51# vdd ALU_1b_2/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1880 gnd ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_2/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1881 ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_2/a_n14_7# ALU_1b_2/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1882 ALU_1b_2/comparator_0/NOR_2/a_n14_7# ALU_1b_2/comparator_0/NOR_2/A vdd ALU_1b_2/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1883 ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/comparator_0/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1884 gnd ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/NOR_3/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1885 ALU_1b_2/comparator_0/NOR_3/out ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/NOR_3/a_n14_7# ALU_1b_2/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1886 ALU_1b_2/comparator_0/NOR_3/a_n14_7# ALU_1b_2/comparator_0/NOR_3/A vdd ALU_1b_2/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1887 ALU_1b_2/comparator_0/NOR_3/out ALU_1b_2/comparator_0/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1888 ALU_1b_2/comparator_0/AND_0/a_78_51# ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1889 ALU_1b_2/comparator_0/NOR_0/A ALU_1b_2/comparator_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1890 vdd ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_0/a_78_51# ALU_1b_2/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1891 ALU_1b_2/comparator_0/AND_0/a_78_51# ALU_1b_2/AND_6/out vdd ALU_1b_2/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1892 ALU_1b_2/comparator_0/AND_0/a_78_8# ALU_1b_2/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1893 ALU_1b_2/comparator_0/NOR_0/A ALU_1b_2/comparator_0/AND_0/a_78_51# vdd ALU_1b_2/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1894 ALU_1b_2/comparator_0/AND_1/a_78_51# ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1895 ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1896 vdd ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/AND_1/a_78_51# ALU_1b_2/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1897 ALU_1b_2/comparator_0/AND_1/a_78_51# ALU_1b_2/AND_6/out vdd ALU_1b_2/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1898 ALU_1b_2/comparator_0/AND_1/a_78_8# ALU_1b_2/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1899 ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/AND_1/a_78_51# vdd ALU_1b_2/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1900 ALU_1b_2/comparator_0/AND_2/a_78_51# ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1901 ALU_1b_2/comparator_0/NOR_1/A ALU_1b_2/comparator_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1902 vdd ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_2/a_78_51# ALU_1b_2/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1903 ALU_1b_2/comparator_0/AND_2/a_78_51# ALU_1b_2/AND_9/out vdd ALU_1b_2/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1904 ALU_1b_2/comparator_0/AND_2/a_78_8# ALU_1b_2/AND_9/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1905 ALU_1b_2/comparator_0/NOR_1/A ALU_1b_2/comparator_0/AND_2/a_78_51# vdd ALU_1b_2/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1906 ALU_1b_2/comparator_0/AND_3/a_78_51# ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1907 ALU_1b_2/comparator_0/NOR_2/A ALU_1b_2/comparator_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1908 vdd ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_3/a_78_51# ALU_1b_2/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1909 ALU_1b_2/comparator_0/AND_3/a_78_51# ALU_1b_2/AND_8/out vdd ALU_1b_2/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1910 ALU_1b_2/comparator_0/AND_3/a_78_8# ALU_1b_2/AND_8/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1911 ALU_1b_2/comparator_0/NOR_2/A ALU_1b_2/comparator_0/AND_3/a_78_51# vdd ALU_1b_2/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1912 ALU_1b_2/comparator_0/AND_5/a_78_51# ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1913 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1914 vdd ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_5/a_78_51# ALU_1b_2/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1915 ALU_1b_2/comparator_0/AND_5/a_78_51# ALU_1b_2/AND_7/out vdd ALU_1b_2/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1916 ALU_1b_2/comparator_0/AND_5/a_78_8# ALU_1b_2/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1917 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_5/a_78_51# vdd ALU_1b_2/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1918 ALU_1b_2/comparator_0/AND_4/a_78_51# ALU_1b_2/AND_8/out ALU_1b_2/comparator_0/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1919 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1920 vdd ALU_1b_2/AND_8/out ALU_1b_2/comparator_0/AND_4/a_78_51# ALU_1b_2/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1921 ALU_1b_2/comparator_0/AND_4/a_78_51# ALU_1b_2/AND_7/out vdd ALU_1b_2/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1922 ALU_1b_2/comparator_0/AND_4/a_78_8# ALU_1b_2/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1923 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_4/a_78_51# vdd ALU_1b_2/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1924 gnd ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1925 ALU_1b_2/comparator_0/NOR_0/out ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/NOR_0/a_n14_7# ALU_1b_2/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1926 ALU_1b_2/comparator_0/NOR_0/a_n14_7# ALU_1b_2/comparator_0/NOR_0/A vdd ALU_1b_2/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1927 ALU_1b_2/comparator_0/NOR_0/out ALU_1b_2/comparator_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1928 gnd ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/comparator_0/NOR_1/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1929 ALU_1b_2/comparator_0/NOR_1/out ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/comparator_0/NOR_1/a_n14_7# ALU_1b_2/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1930 ALU_1b_2/comparator_0/NOR_1/a_n14_7# ALU_1b_2/comparator_0/NOR_1/A vdd ALU_1b_2/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1931 ALU_1b_2/comparator_0/NOR_1/out ALU_1b_2/comparator_0/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1932 vdd ALU_1b_2/comparator_0/NOR_1/out ALU_1b_2/AND_10/B ALU_1b_2/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1933 gnd ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_5/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1934 gnd ALU_1b_2/comparator_0/NOR_0/out ALU_1b_2/comparator_0/NOR_1/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1935 vdd ALU_1b_2/comparator_0/NOR_0/out ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1936 gnd ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/AND_11/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1937 vdd ALU_1b_2/comparator_0/NOR_3/out ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=9 ps=5
M1938 gnd ALU_1b_2/comparator_0/NOR_3/out ALU_1b_2/comparator_0/NOR_2/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1939 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1940 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/AND_7/out vdd ALU_1b_2/comparator_0/w_n39_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1941 gnd ALU_1b_2/comparator_0/NOR_1/out ALU_1b_2/AND_10/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1942 vdd ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/AND_11/B ALU_1b_2/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1943 vdd ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/w_n74_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=1 ps=1
M1944 ALU_1b_2/AND_19/A ALU_1b_2/NOT_1/in vdd ALU_1b_2/NOT_1/w_n36_43# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1945 ALU_1b_2/AND_19/A ALU_1b_2/NOT_1/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1946 ALU_1b_2/AND_3/A A1 vdd ALU_1b_2/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1947 ALU_1b_2/AND_3/A A1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1948 ALU_1b_2/NOR_2/A ALU_1b_2/NOT_2/in vdd ALU_1b_2/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1949 ALU_1b_2/NOR_2/A ALU_1b_2/NOT_2/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1950 ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/decoder_0/AND_1/B ALU_1b_2/decoder_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1951 ALU_1b_2/AND_2/B ALU_1b_2/decoder_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1952 vdd ALU_1b_2/decoder_0/AND_1/B ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1953 ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/decoder_0/AND_2/B vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1954 ALU_1b_2/decoder_0/AND_0/a_78_8# ALU_1b_2/decoder_0/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1955 ALU_1b_2/AND_2/B ALU_1b_2/decoder_0/AND_0/a_78_51# vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1956 ALU_1b_2/decoder_0/AND_1/a_78_51# ALU_1b_2/decoder_0/AND_1/B ALU_1b_2/decoder_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1957 ALU_1b_2/AND_9/A ALU_1b_2/decoder_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1958 vdd ALU_1b_2/decoder_0/AND_1/B ALU_1b_2/decoder_0/AND_1/a_78_51# ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1959 ALU_1b_2/decoder_0/AND_1/a_78_51# S1 vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 ALU_1b_2/decoder_0/AND_1/a_78_8# S1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1961 ALU_1b_2/AND_9/A ALU_1b_2/decoder_0/AND_1/a_78_51# vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1962 ALU_1b_2/decoder_0/AND_2/a_78_51# ALU_1b_2/decoder_0/AND_2/B ALU_1b_2/decoder_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1963 ALU_1b_2/AND_5/B ALU_1b_2/decoder_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1964 vdd ALU_1b_2/decoder_0/AND_2/B ALU_1b_2/decoder_0/AND_2/a_78_51# ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1965 ALU_1b_2/decoder_0/AND_2/a_78_51# S0 vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1966 ALU_1b_2/decoder_0/AND_2/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1967 ALU_1b_2/AND_5/B ALU_1b_2/decoder_0/AND_2/a_78_51# vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1968 ALU_1b_2/decoder_0/AND_3/a_78_51# S1 ALU_1b_2/decoder_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M1969 ALU_1b_2/AND_15/A ALU_1b_2/decoder_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1970 vdd S1 ALU_1b_2/decoder_0/AND_3/a_78_51# ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1971 ALU_1b_2/decoder_0/AND_3/a_78_51# S0 vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1972 ALU_1b_2/decoder_0/AND_3/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1973 ALU_1b_2/AND_15/A ALU_1b_2/decoder_0/AND_3/a_78_51# vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1974 ALU_1b_2/decoder_0/AND_2/B S1 vdd ALU_1b_2/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1975 ALU_1b_2/decoder_0/AND_2/B S1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1976 ALU_1b_2/decoder_0/AND_1/B S0 vdd ALU_1b_2/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1977 ALU_1b_2/decoder_0/AND_1/B S0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1978 ALU_1b_2/NOR_2/B ALU_1b_2/NOT_3/in vdd ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1979 ALU_1b_2/NOR_2/B ALU_1b_2/NOT_3/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1980 gnd ALU_1b_2/NOR_0/B ALU_1b_2/NOT_2/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1981 ALU_1b_2/NOT_2/in ALU_1b_2/NOR_0/B ALU_1b_2/NOR_0/a_n14_7# ALU_1b_2/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1982 ALU_1b_2/NOR_0/a_n14_7# ALU_1b_2/NOR_0/A vdd ALU_1b_2/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1983 ALU_1b_2/NOT_2/in ALU_1b_2/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1984 F1 ALU_1b_2/NOT_4/in vdd ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1985 F1 ALU_1b_2/NOT_4/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1986 gnd ALU_1b_2/NOR_1/B ALU_1b_2/NOT_3/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1987 ALU_1b_2/NOT_3/in ALU_1b_2/NOR_1/B ALU_1b_2/NOR_1/a_n14_7# ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1988 ALU_1b_2/NOR_1/a_n14_7# ALU_1b_2/NOR_1/A vdd ALU_1b_2/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1989 ALU_1b_2/NOT_3/in ALU_1b_2/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1990 gnd ALU_1b_3/NOR_2/B ALU_1b_3/NOT_4/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1991 ALU_1b_3/NOT_4/in ALU_1b_3/NOR_2/B ALU_1b_3/NOR_2/a_n14_7# ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1992 ALU_1b_3/NOR_2/a_n14_7# ALU_1b_3/NOR_2/A vdd ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1993 ALU_1b_3/NOT_4/in ALU_1b_3/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1994 ALU_1b_3/NOR_4/B ALU_1b_3/NOT_5/in vdd ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1995 ALU_1b_3/NOR_4/B ALU_1b_3/NOT_5/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1996 ALU_1b_1/C0 ALU_1b_3/NOT_6/in vdd ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1997 ALU_1b_1/C0 ALU_1b_3/NOT_6/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M1998 gnd ALU_1b_3/NOR_3/B ALU_1b_3/NOT_5/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1999 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_3/B ALU_1b_3/NOR_3/a_n14_7# ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2000 ALU_1b_3/NOR_3/a_n14_7# ALU_1b_3/NOR_3/A vdd ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2001 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2002 gnd ALU_1b_3/NOR_4/B ALU_1b_3/NOT_6/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2003 ALU_1b_3/NOT_6/in ALU_1b_3/NOR_4/B ALU_1b_3/NOR_4/a_n14_7# ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2004 ALU_1b_3/NOR_4/a_n14_7# ALU_1b_3/NOR_4/A vdd ALU_1b_3/NOR_4/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2005 ALU_1b_3/NOT_6/in ALU_1b_3/NOR_4/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2006 ALU_1b_3/AND_0/a_78_51# A2 ALU_1b_3/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2007 ALU_1b_3/AND_0/out ALU_1b_3/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2008 vdd A2 ALU_1b_3/AND_0/a_78_51# ALU_1b_3/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2009 ALU_1b_3/AND_0/a_78_51# ALU_1b_3/AND_2/B vdd ALU_1b_3/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2010 ALU_1b_3/AND_0/a_78_8# ALU_1b_3/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2011 ALU_1b_3/AND_0/out ALU_1b_3/AND_0/a_78_51# vdd ALU_1b_3/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2012 ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2013 ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out ALU_1b_3/full_adder_0/half_adder_1/A vdd ALU_1b_3/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M2014 vdd ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out ALU_1b_3/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2015 ALU_1b_3/full_adder_0/half_adder_1/NAND_0/a_n7_n34# ALU_1b_3/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2016 ALU_1b_3/AND_16/A ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2017 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_0/half_adder_1/A vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2018 ALU_1b_3/AND_16/A ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2019 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_3/AND_1/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2020 gnd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2021 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2022 vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2023 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/AND_16/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2024 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_74# ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_16/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2025 gnd ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2026 vdd ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2027 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_0/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2028 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out vdd ALU_1b_3/full_adder_0/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2029 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2030 ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2031 ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out ALU_1b_3/AND_0/out vdd ALU_1b_3/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M2032 vdd ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out ALU_1b_3/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2033 ALU_1b_3/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_3/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2034 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2035 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_3/AND_0/out vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2036 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2037 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# ALU_1b_3/AND_2/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2038 gnd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2039 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2040 vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2041 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_3/full_adder_0/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2042 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2043 gnd ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2044 vdd ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2045 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_3/AND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2046 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out vdd ALU_1b_3/full_adder_0/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2047 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2048 gnd ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2049 ALU_1b_3/full_adder_0/NOR_0/out ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/NOR_0/a_n14_7# ALU_1b_3/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2050 ALU_1b_3/full_adder_0/NOR_0/a_n14_7# ALU_1b_3/full_adder_0/NOR_0/A vdd ALU_1b_3/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2051 ALU_1b_3/full_adder_0/NOR_0/out ALU_1b_3/full_adder_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2052 ALU_1b_3/AND_17/A ALU_1b_3/full_adder_0/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2053 ALU_1b_3/AND_17/A ALU_1b_3/full_adder_0/NOR_0/out vdd ALU_1b_3/full_adder_0/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2054 ALU_1b_3/AND_1/a_78_51# ALU_1b_3/AND_2/B ALU_1b_3/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2055 ALU_1b_3/AND_1/out ALU_1b_3/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2056 vdd ALU_1b_3/AND_2/B ALU_1b_3/AND_1/a_78_51# ALU_1b_3/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2057 ALU_1b_3/AND_1/a_78_51# ALU_1b_3/C0 vdd ALU_1b_3/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2058 ALU_1b_3/AND_1/a_78_8# ALU_1b_3/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2059 ALU_1b_3/AND_1/out ALU_1b_3/AND_1/a_78_51# vdd ALU_1b_3/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2060 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2061 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/full_adder_1/half_adder_1/A vdd ALU_1b_3/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M2062 vdd ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2063 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/a_n7_n34# ALU_1b_3/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2064 ALU_1b_3/NOT_1/in ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2065 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_1/half_adder_1/A vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2066 ALU_1b_3/NOT_1/in ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2067 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_3/AND_5/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2068 gnd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2069 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2070 vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2071 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_3/NOT_1/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2072 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/NOT_1/in ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2073 gnd ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2074 vdd ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2075 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_1/half_adder_1/A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2076 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out vdd ALU_1b_3/full_adder_1/half_adder_1/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2077 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2078 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/NAND_0/a_n7_n34# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2079 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/AND_3/out vdd ALU_1b_3/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M2080 vdd ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2081 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_3/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2082 ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/AND_3/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2083 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_3/AND_3/out vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2084 ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M2085 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_3/AND_4/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2086 gnd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2087 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2088 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2089 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_3/full_adder_1/half_adder_1/A Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2090 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_3/AND_3/out ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2091 gnd ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2092 vdd ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2093 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_3/AND_3/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2094 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out vdd ALU_1b_3/full_adder_1/half_adder_0/w_36_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2095 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2096 gnd ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2097 ALU_1b_3/full_adder_1/NOR_0/out ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/NOR_0/a_n14_7# ALU_1b_3/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2098 ALU_1b_3/full_adder_1/NOR_0/a_n14_7# ALU_1b_3/full_adder_1/NOR_0/A vdd ALU_1b_3/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2099 ALU_1b_3/full_adder_1/NOR_0/out ALU_1b_3/full_adder_1/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2100 ALU_1b_3/AND_18/A ALU_1b_3/full_adder_1/NOR_0/out gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2101 ALU_1b_3/AND_18/A ALU_1b_3/full_adder_1/NOR_0/out vdd ALU_1b_3/full_adder_1/w_448_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2102 ALU_1b_3/AND_2/a_78_51# ALU_1b_3/AND_2/B ALU_1b_3/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2103 ALU_1b_3/AND_2/out ALU_1b_3/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2104 vdd ALU_1b_3/AND_2/B ALU_1b_3/AND_2/a_78_51# ALU_1b_3/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2105 ALU_1b_3/AND_2/a_78_51# B2 vdd ALU_1b_3/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2106 ALU_1b_3/AND_2/a_78_8# B2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2107 ALU_1b_3/AND_2/out ALU_1b_3/AND_2/a_78_51# vdd ALU_1b_3/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2108 ALU_1b_3/AND_3/a_78_51# ALU_1b_3/AND_5/B ALU_1b_3/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2109 ALU_1b_3/AND_3/out ALU_1b_3/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2110 vdd ALU_1b_3/AND_5/B ALU_1b_3/AND_3/a_78_51# ALU_1b_3/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2111 ALU_1b_3/AND_3/a_78_51# ALU_1b_3/AND_3/A vdd ALU_1b_3/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2112 ALU_1b_3/AND_3/a_78_8# ALU_1b_3/AND_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2113 ALU_1b_3/AND_3/out ALU_1b_3/AND_3/a_78_51# vdd ALU_1b_3/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2114 ALU_1b_3/AND_5/a_78_51# ALU_1b_3/AND_5/B ALU_1b_3/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2115 ALU_1b_3/AND_5/out ALU_1b_3/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2116 vdd ALU_1b_3/AND_5/B ALU_1b_3/AND_5/a_78_51# ALU_1b_3/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2117 ALU_1b_3/AND_5/a_78_51# ALU_1b_3/C0 vdd ALU_1b_3/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2118 ALU_1b_3/AND_5/a_78_8# ALU_1b_3/C0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2119 ALU_1b_3/AND_5/out ALU_1b_3/AND_5/a_78_51# vdd ALU_1b_3/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2120 ALU_1b_3/AND_4/a_78_51# ALU_1b_3/AND_5/B ALU_1b_3/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2121 ALU_1b_3/AND_4/out ALU_1b_3/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2122 vdd ALU_1b_3/AND_5/B ALU_1b_3/AND_4/a_78_51# ALU_1b_3/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2123 ALU_1b_3/AND_4/a_78_51# B2 vdd ALU_1b_3/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2124 ALU_1b_3/AND_4/a_78_8# B2 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2125 ALU_1b_3/AND_4/out ALU_1b_3/AND_4/a_78_51# vdd ALU_1b_3/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2126 ALU_1b_3/AND_10/a_78_51# ALU_1b_3/AND_10/B ALU_1b_3/AND_10/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2127 ALU_1b_3/NOR_1/A ALU_1b_3/AND_10/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2128 vdd ALU_1b_3/AND_10/B ALU_1b_3/AND_10/a_78_51# ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2129 ALU_1b_3/AND_10/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2130 ALU_1b_3/AND_10/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2131 ALU_1b_3/NOR_1/A ALU_1b_3/AND_10/a_78_51# vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2132 ALU_1b_3/AND_11/a_78_51# ALU_1b_3/AND_11/B ALU_1b_3/AND_11/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2133 ALU_1b_3/NOR_4/A ALU_1b_3/AND_11/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2134 vdd ALU_1b_3/AND_11/B ALU_1b_3/AND_11/a_78_51# ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2135 ALU_1b_3/AND_11/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2136 ALU_1b_3/AND_11/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2137 ALU_1b_3/NOR_4/A ALU_1b_3/AND_11/a_78_51# vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2138 ALU_1b_3/AND_6/a_78_51# A2 ALU_1b_3/AND_6/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2139 ALU_1b_3/AND_6/out ALU_1b_3/AND_6/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2140 vdd A2 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2141 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2142 ALU_1b_3/AND_6/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2143 ALU_1b_3/AND_6/out ALU_1b_3/AND_6/a_78_51# vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2144 ALU_1b_3/AND_7/a_78_51# B2 ALU_1b_3/AND_7/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2145 ALU_1b_3/AND_7/out ALU_1b_3/AND_7/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2146 vdd B2 ALU_1b_3/AND_7/a_78_51# ALU_1b_3/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2147 ALU_1b_3/AND_7/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2148 ALU_1b_3/AND_7/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2149 ALU_1b_3/AND_7/out ALU_1b_3/AND_7/a_78_51# vdd ALU_1b_3/AND_7/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2150 ALU_1b_3/AND_12/a_78_51# A2 ALU_1b_3/AND_12/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2151 ALU_1b_3/AND_14/B ALU_1b_3/AND_12/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2152 vdd A2 ALU_1b_3/AND_12/a_78_51# ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2153 ALU_1b_3/AND_12/a_78_51# ALU_1b_3/AND_15/A vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2154 ALU_1b_3/AND_12/a_78_8# ALU_1b_3/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2155 ALU_1b_3/AND_14/B ALU_1b_3/AND_12/a_78_51# vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2156 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/C0 ALU_1b_3/AND_8/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2157 ALU_1b_3/AND_8/out ALU_1b_3/AND_8/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2158 vdd ALU_1b_3/C0 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2159 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2160 ALU_1b_3/AND_8/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2161 ALU_1b_3/AND_8/out ALU_1b_3/AND_8/a_78_51# vdd ALU_1b_3/AND_8/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2162 ALU_1b_3/AND_13/a_78_51# B2 ALU_1b_3/AND_13/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2163 ALU_1b_3/AND_14/A ALU_1b_3/AND_13/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2164 vdd B2 ALU_1b_3/AND_13/a_78_51# ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2165 ALU_1b_3/AND_13/a_78_51# ALU_1b_3/AND_15/A vdd ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2166 ALU_1b_3/AND_13/a_78_8# ALU_1b_3/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2167 ALU_1b_3/AND_14/A ALU_1b_3/AND_13/a_78_51# vdd ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2168 ALU_1b_3/AND_9/a_78_51# F1 ALU_1b_3/AND_9/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2169 ALU_1b_3/AND_9/out ALU_1b_3/AND_9/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2170 vdd F1 ALU_1b_3/AND_9/a_78_51# ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2171 ALU_1b_3/AND_9/a_78_51# ALU_1b_3/AND_9/A vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2172 ALU_1b_3/AND_9/a_78_8# ALU_1b_3/AND_9/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2173 ALU_1b_3/AND_9/out ALU_1b_3/AND_9/a_78_51# vdd ALU_1b_3/AND_9/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2174 ALU_1b_3/AND_14/a_78_51# ALU_1b_3/AND_14/B ALU_1b_3/AND_14/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2175 ALU_1b_3/AND_15/B ALU_1b_3/AND_14/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2176 vdd ALU_1b_3/AND_14/B ALU_1b_3/AND_14/a_78_51# ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2177 ALU_1b_3/AND_14/a_78_51# ALU_1b_3/AND_14/A vdd ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2178 ALU_1b_3/AND_14/a_78_8# ALU_1b_3/AND_14/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2179 ALU_1b_3/AND_15/B ALU_1b_3/AND_14/a_78_51# vdd ALU_1b_3/AND_14/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2180 ALU_1b_3/AND_15/a_78_51# ALU_1b_3/AND_15/B ALU_1b_3/AND_15/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2181 ALU_1b_3/NOR_1/B ALU_1b_3/AND_15/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2182 vdd ALU_1b_3/AND_15/B ALU_1b_3/AND_15/a_78_51# ALU_1b_3/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2183 ALU_1b_3/AND_15/a_78_51# ALU_1b_3/AND_15/A vdd ALU_1b_3/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2184 ALU_1b_3/AND_15/a_78_8# ALU_1b_3/AND_15/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2185 ALU_1b_3/NOR_1/B ALU_1b_3/AND_15/a_78_51# vdd ALU_1b_3/AND_15/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2186 ALU_1b_3/AND_16/a_78_51# ALU_1b_3/AND_2/B ALU_1b_3/AND_16/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2187 ALU_1b_3/NOR_0/B ALU_1b_3/AND_16/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2188 vdd ALU_1b_3/AND_2/B ALU_1b_3/AND_16/a_78_51# ALU_1b_3/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2189 ALU_1b_3/AND_16/a_78_51# ALU_1b_3/AND_16/A vdd ALU_1b_3/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2190 ALU_1b_3/AND_16/a_78_8# ALU_1b_3/AND_16/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2191 ALU_1b_3/NOR_0/B ALU_1b_3/AND_16/a_78_51# vdd ALU_1b_3/AND_16/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2192 ALU_1b_3/AND_17/a_78_51# ALU_1b_3/AND_2/B ALU_1b_3/AND_17/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2193 ALU_1b_3/NOR_3/B ALU_1b_3/AND_17/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2194 vdd ALU_1b_3/AND_2/B ALU_1b_3/AND_17/a_78_51# ALU_1b_3/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2195 ALU_1b_3/AND_17/a_78_51# ALU_1b_3/AND_17/A vdd ALU_1b_3/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2196 ALU_1b_3/AND_17/a_78_8# ALU_1b_3/AND_17/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2197 ALU_1b_3/NOR_3/B ALU_1b_3/AND_17/a_78_51# vdd ALU_1b_3/AND_17/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2198 ALU_1b_3/AND_19/a_78_51# ALU_1b_3/AND_5/B ALU_1b_3/AND_19/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2199 ALU_1b_3/NOR_0/A ALU_1b_3/AND_19/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2200 vdd ALU_1b_3/AND_5/B ALU_1b_3/AND_19/a_78_51# ALU_1b_3/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2201 ALU_1b_3/AND_19/a_78_51# ALU_1b_3/AND_19/A vdd ALU_1b_3/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2202 ALU_1b_3/AND_19/a_78_8# ALU_1b_3/AND_19/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2203 ALU_1b_3/NOR_0/A ALU_1b_3/AND_19/a_78_51# vdd ALU_1b_3/AND_19/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2204 ALU_1b_3/AND_18/a_78_51# ALU_1b_3/AND_5/B ALU_1b_3/AND_18/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2205 ALU_1b_3/NOR_3/A ALU_1b_3/AND_18/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2206 vdd ALU_1b_3/AND_5/B ALU_1b_3/AND_18/a_78_51# ALU_1b_3/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2207 ALU_1b_3/AND_18/a_78_51# ALU_1b_3/AND_18/A vdd ALU_1b_3/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2208 ALU_1b_3/AND_18/a_78_8# ALU_1b_3/AND_18/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2209 ALU_1b_3/NOR_3/A ALU_1b_3/AND_18/a_78_51# vdd ALU_1b_3/AND_18/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2210 gnd ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_2/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2211 ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_2/a_n14_7# ALU_1b_3/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2212 ALU_1b_3/comparator_0/NOR_2/a_n14_7# ALU_1b_3/comparator_0/NOR_2/A vdd ALU_1b_3/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2213 ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/comparator_0/NOR_2/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2214 gnd ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/NOR_3/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2215 ALU_1b_3/comparator_0/NOR_3/out ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/NOR_3/a_n14_7# ALU_1b_3/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2216 ALU_1b_3/comparator_0/NOR_3/a_n14_7# ALU_1b_3/comparator_0/NOR_3/A vdd ALU_1b_3/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2217 ALU_1b_3/comparator_0/NOR_3/out ALU_1b_3/comparator_0/NOR_3/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2218 ALU_1b_3/comparator_0/AND_0/a_78_51# ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2219 ALU_1b_3/comparator_0/NOR_0/A ALU_1b_3/comparator_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2220 vdd ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_0/a_78_51# ALU_1b_3/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2221 ALU_1b_3/comparator_0/AND_0/a_78_51# ALU_1b_3/AND_6/out vdd ALU_1b_3/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2222 ALU_1b_3/comparator_0/AND_0/a_78_8# ALU_1b_3/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2223 ALU_1b_3/comparator_0/NOR_0/A ALU_1b_3/comparator_0/AND_0/a_78_51# vdd ALU_1b_3/comparator_0/AND_0/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2224 ALU_1b_3/comparator_0/AND_1/a_78_51# ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2225 ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2226 vdd ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/AND_1/a_78_51# ALU_1b_3/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2227 ALU_1b_3/comparator_0/AND_1/a_78_51# ALU_1b_3/AND_6/out vdd ALU_1b_3/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2228 ALU_1b_3/comparator_0/AND_1/a_78_8# ALU_1b_3/AND_6/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2229 ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/AND_1/a_78_51# vdd ALU_1b_3/comparator_0/AND_1/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2230 ALU_1b_3/comparator_0/AND_2/a_78_51# ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2231 ALU_1b_3/comparator_0/NOR_1/A ALU_1b_3/comparator_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2232 vdd ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_2/a_78_51# ALU_1b_3/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2233 ALU_1b_3/comparator_0/AND_2/a_78_51# ALU_1b_3/AND_9/out vdd ALU_1b_3/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2234 ALU_1b_3/comparator_0/AND_2/a_78_8# ALU_1b_3/AND_9/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2235 ALU_1b_3/comparator_0/NOR_1/A ALU_1b_3/comparator_0/AND_2/a_78_51# vdd ALU_1b_3/comparator_0/AND_2/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2236 ALU_1b_3/comparator_0/AND_3/a_78_51# ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2237 ALU_1b_3/comparator_0/NOR_2/A ALU_1b_3/comparator_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2238 vdd ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_3/a_78_51# ALU_1b_3/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2239 ALU_1b_3/comparator_0/AND_3/a_78_51# ALU_1b_3/AND_8/out vdd ALU_1b_3/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2240 ALU_1b_3/comparator_0/AND_3/a_78_8# ALU_1b_3/AND_8/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2241 ALU_1b_3/comparator_0/NOR_2/A ALU_1b_3/comparator_0/AND_3/a_78_51# vdd ALU_1b_3/comparator_0/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2242 ALU_1b_3/comparator_0/AND_5/a_78_51# ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_5/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2243 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_5/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2244 vdd ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_5/a_78_51# ALU_1b_3/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2245 ALU_1b_3/comparator_0/AND_5/a_78_51# ALU_1b_3/AND_7/out vdd ALU_1b_3/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2246 ALU_1b_3/comparator_0/AND_5/a_78_8# ALU_1b_3/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2247 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_5/a_78_51# vdd ALU_1b_3/comparator_0/AND_5/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2248 ALU_1b_3/comparator_0/AND_4/a_78_51# ALU_1b_3/AND_8/out ALU_1b_3/comparator_0/AND_4/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2249 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_4/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2250 vdd ALU_1b_3/AND_8/out ALU_1b_3/comparator_0/AND_4/a_78_51# ALU_1b_3/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2251 ALU_1b_3/comparator_0/AND_4/a_78_51# ALU_1b_3/AND_7/out vdd ALU_1b_3/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2252 ALU_1b_3/comparator_0/AND_4/a_78_8# ALU_1b_3/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2253 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_4/a_78_51# vdd ALU_1b_3/comparator_0/AND_4/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2254 gnd ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/NOR_0/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2255 ALU_1b_3/comparator_0/NOR_0/out ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/NOR_0/a_n14_7# ALU_1b_3/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2256 ALU_1b_3/comparator_0/NOR_0/a_n14_7# ALU_1b_3/comparator_0/NOR_0/A vdd ALU_1b_3/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2257 ALU_1b_3/comparator_0/NOR_0/out ALU_1b_3/comparator_0/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2258 gnd ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/comparator_0/NOR_1/out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2259 ALU_1b_3/comparator_0/NOR_1/out ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/comparator_0/NOR_1/a_n14_7# ALU_1b_3/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2260 ALU_1b_3/comparator_0/NOR_1/a_n14_7# ALU_1b_3/comparator_0/NOR_1/A vdd ALU_1b_3/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2261 ALU_1b_3/comparator_0/NOR_1/out ALU_1b_3/comparator_0/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2262 vdd ALU_1b_3/comparator_0/NOR_1/out ALU_1b_3/AND_10/B ALU_1b_3/comparator_0/w_113_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2263 gnd ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_5/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2264 gnd ALU_1b_3/comparator_0/NOR_0/out ALU_1b_3/comparator_0/NOR_1/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2265 vdd ALU_1b_3/comparator_0/NOR_0/out ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/comparator_0/w_88_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2266 gnd ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/AND_11/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2267 vdd ALU_1b_3/comparator_0/NOR_3/out ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/w_n195_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=9 ps=5
M2268 gnd ALU_1b_3/comparator_0/NOR_3/out ALU_1b_3/comparator_0/NOR_2/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2269 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/AND_7/out gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2270 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/AND_7/out vdd ALU_1b_3/comparator_0/w_n39_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2271 gnd ALU_1b_3/comparator_0/NOR_1/out ALU_1b_3/AND_10/B Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2272 vdd ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/AND_11/B ALU_1b_3/comparator_0/w_n220_n67# CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M2273 vdd ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/w_n74_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=1 ps=1
M2274 ALU_1b_3/AND_19/A ALU_1b_3/NOT_1/in vdd ALU_1b_3/NOT_1/w_n36_43# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2275 ALU_1b_3/AND_19/A ALU_1b_3/NOT_1/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2276 ALU_1b_3/AND_3/A A2 vdd ALU_1b_3/AND_3/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2277 ALU_1b_3/AND_3/A A2 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2278 ALU_1b_3/NOR_2/A ALU_1b_3/NOT_2/in vdd ALU_1b_3/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2279 ALU_1b_3/NOR_2/A ALU_1b_3/NOT_2/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2280 ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/decoder_0/AND_1/B ALU_1b_3/decoder_0/AND_0/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2281 ALU_1b_3/AND_2/B ALU_1b_3/decoder_0/AND_0/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2282 vdd ALU_1b_3/decoder_0/AND_1/B ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2283 ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/decoder_0/AND_2/B vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2284 ALU_1b_3/decoder_0/AND_0/a_78_8# ALU_1b_3/decoder_0/AND_2/B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2285 ALU_1b_3/AND_2/B ALU_1b_3/decoder_0/AND_0/a_78_51# vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2286 ALU_1b_3/decoder_0/AND_1/a_78_51# ALU_1b_3/decoder_0/AND_1/B ALU_1b_3/decoder_0/AND_1/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2287 ALU_1b_3/AND_9/A ALU_1b_3/decoder_0/AND_1/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2288 vdd ALU_1b_3/decoder_0/AND_1/B ALU_1b_3/decoder_0/AND_1/a_78_51# ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2289 ALU_1b_3/decoder_0/AND_1/a_78_51# S1 vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2290 ALU_1b_3/decoder_0/AND_1/a_78_8# S1 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2291 ALU_1b_3/AND_9/A ALU_1b_3/decoder_0/AND_1/a_78_51# vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2292 ALU_1b_3/decoder_0/AND_2/a_78_51# ALU_1b_3/decoder_0/AND_2/B ALU_1b_3/decoder_0/AND_2/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2293 ALU_1b_3/AND_5/B ALU_1b_3/decoder_0/AND_2/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2294 vdd ALU_1b_3/decoder_0/AND_2/B ALU_1b_3/decoder_0/AND_2/a_78_51# ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2295 ALU_1b_3/decoder_0/AND_2/a_78_51# S0 vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2296 ALU_1b_3/decoder_0/AND_2/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2297 ALU_1b_3/AND_5/B ALU_1b_3/decoder_0/AND_2/a_78_51# vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2298 ALU_1b_3/decoder_0/AND_3/a_78_51# S1 ALU_1b_3/decoder_0/AND_3/a_78_8# Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=32 ps=24
M2299 ALU_1b_3/AND_15/A ALU_1b_3/decoder_0/AND_3/a_78_51# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2300 vdd S1 ALU_1b_3/decoder_0/AND_3/a_78_51# ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M2301 ALU_1b_3/decoder_0/AND_3/a_78_51# S0 vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2302 ALU_1b_3/decoder_0/AND_3/a_78_8# S0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2303 ALU_1b_3/AND_15/A ALU_1b_3/decoder_0/AND_3/a_78_51# vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M2304 ALU_1b_3/decoder_0/AND_2/B S1 vdd ALU_1b_3/AND_6/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2305 ALU_1b_3/decoder_0/AND_2/B S1 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2306 ALU_1b_3/decoder_0/AND_1/B S0 vdd ALU_1b_3/AND_12/w_64_45# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2307 ALU_1b_3/decoder_0/AND_1/B S0 gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2308 ALU_1b_3/NOR_2/B ALU_1b_3/NOT_3/in vdd ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2309 ALU_1b_3/NOR_2/B ALU_1b_3/NOT_3/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2310 gnd ALU_1b_3/NOR_0/B ALU_1b_3/NOT_2/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2311 ALU_1b_3/NOT_2/in ALU_1b_3/NOR_0/B ALU_1b_3/NOR_0/a_n14_7# ALU_1b_3/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2312 ALU_1b_3/NOR_0/a_n14_7# ALU_1b_3/NOR_0/A vdd ALU_1b_3/NOR_0/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2313 ALU_1b_3/NOT_2/in ALU_1b_3/NOR_0/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2314 F2 ALU_1b_3/NOT_4/in vdd ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2315 F2 ALU_1b_3/NOT_4/in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
M2316 gnd ALU_1b_3/NOR_1/B ALU_1b_3/NOT_3/in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M2317 ALU_1b_3/NOT_3/in ALU_1b_3/NOR_1/B ALU_1b_3/NOR_1/a_n14_7# ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M2318 ALU_1b_3/NOR_1/a_n14_7# ALU_1b_3/NOR_1/A vdd ALU_1b_3/NOR_2/w_n27_1# CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M2319 ALU_1b_3/NOT_3/in ALU_1b_3/NOR_1/A gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A1 ALU_1b_2/AND_3/A 0.03fF
C1 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_2/out 0.27fF
C2 vdd ALU_1b_3/full_adder_1/w_448_45# 0.12fF
C3 ALU_1b_0/AND_14/B B0 0.23fF
C4 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_1/out 0.72fF
C5 ALU_1b_2/AND_10/a_78_51# ALU_1b_2/AND_10/B 0.38fF
C6 ALU_1b_3/AND_15/a_78_51# ALU_1b_3/NOR_1/B 0.05fF
C7 ALU_1b_0/AND_5/a_78_51# ALU_1b_0/AND_5/B 0.19fF
C8 ALU_1b_0/decoder_0/AND_2/B ALU_1b_0/AND_12/w_64_45# 0.06fF
C9 ALU_1b_0/NOR_4/A ALU_1b_0/NOR_4/B 0.35fF
C10 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C11 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_6/out 0.05fF
C12 gnd ALU_1b_3/AND_0/a_78_51# 0.07fF
C13 S1 ALU_1b_1/decoder_0/AND_2/B 0.07fF
C14 ALU_1b_1/AND_9/A B3 0.28fF
C15 ALU_1b_1/NOR_0/A gnd 0.17fF
C16 vdd ALU_1b_3/AND_18/w_64_45# 0.15fF
C17 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/NOT_1/in 0.23fF
C18 ALU_1b_3/AND_5/w_64_45# ALU_1b_3/AND_5/B 0.06fF
C19 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_1/NOR_0/A 0.06fF
C20 ALU_1b_0/AND_4/out gnd 0.07fF
C21 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C22 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/NOR_0/B 0.09fF
C23 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C24 gnd ALU_1b_3/AND_18/a_78_51# 0.07fF
C25 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_2/AND_16/A 0.13fF
C26 vdd ALU_1b_2/comparator_0/NOR_1/A 0.03fF
C27 ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C28 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C29 ALU_1b_1/AND_5/out vdd 0.35fF
C30 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/A 0.16fF
C31 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.00fF
C32 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/NOR_0/A 0.10fF
C33 gnd ALU_1b_3/AND_2/B 0.48fF
C34 ALU_1b_0/full_adder_1/w_448_45# ALU_1b_0/AND_18/A 0.03fF
C35 ALU_1b_1/comparator_0/w_n220_n67# ALU_1b_1/comparator_0/NOR_2/A 0.06fF
C36 A3 ALU_1b_1/AND_12/a_78_51# 0.19fF
C37 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C38 ALU_1b_3/AND_4/out F1 0.01fF
C39 ALU_1b_0/AND_19/w_64_45# ALU_1b_0/NOR_0/A 0.03fF
C40 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/AND_1/out 0.70fF
C41 ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/AND_1/a_78_51# 0.20fF
C42 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_2/a_78_51# 0.19fF
C43 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_5/B 0.17fF
C44 ALU_1b_0/AND_14/A gnd 0.07fF
C45 vdd ALU_1b_2/AND_8/out 0.66fF
C46 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_9/a_78_51# 0.09fF
C47 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C48 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/AND_5/out 0.20fF
C49 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/AND_3/out 0.00fF
C50 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/AND_16/A 0.06fF
C51 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_5/B 0.05fF
C52 ALU_1b_2/decoder_0/AND_2/B ALU_1b_2/decoder_0/AND_1/B 0.59fF
C53 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/NOR_0/B 0.38fF
C54 ALU_1b_0/comparator_0/NOR_1/B vdd 0.30fF
C55 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_1/A 0.13fF
C56 ALU_1b_0/AND_15/B vdd 0.09fF
C57 ALU_1b_3/full_adder_1/half_adder_1/w_36_45# ALU_1b_3/AND_5/out 0.29fF
C58 ALU_1b_1/NOT_2/in ALU_1b_1/NOR_2/A 0.03fF
C59 ALU_1b_1/comparator_0/NOR_2/B gnd 0.07fF
C60 ALU_1b_2/AND_6/out ALU_1b_2/AND_7/out 0.13fF
C61 ALU_1b_0/comparator_0/AND_3/w_64_45# ALU_1b_0/comparator_0/AND_3/a_78_51# 0.09fF
C62 ALU_1b_0/comparator_0/NOR_1/out gnd 0.07fF
C63 ALU_1b_0/AND_9/out ALU_1b_0/AND_7/out 0.02fF
C64 vdd ALU_1b_3/AND_10/a_78_51# 0.06fF
C65 ALU_1b_0/AND_12/a_78_51# ALU_1b_0/AND_15/A 0.05fF
C66 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/AND_3/out 0.23fF
C67 vdd ALU_1b_2/AND_15/a_78_51# 0.06fF
C68 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_3/B 0.15fF
C69 ALU_1b_1/NOT_1/in ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.13fF
C70 gnd ALU_1b_3/comparator_0/NOR_3/A 0.21fF
C71 ALU_1b_1/NOR_0/A ALU_1b_1/NOR_3/A 0.01fF
C72 ALU_1b_3/NOT_3/in ALU_1b_3/NOR_2/w_n27_1# 0.11fF
C73 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/AND_1/out 0.08fF
C74 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_7/out 0.20fF
C75 A2 ALU_1b_3/AND_8/out 0.11fF
C76 ALU_1b_1/AND_9/a_78_51# ALU_1b_1/AND_9/out 0.05fF
C77 ALU_1b_1/AND_7/a_78_51# ALU_1b_1/AND_8/out 0.10fF
C78 A3 vdd 0.21fF
C79 ALU_1b_1/comparator_0/w_113_n67# ALU_1b_1/AND_10/B 0.03fF
C80 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_1/full_adder_0/half_adder_1/A 0.03fF
C81 ALU_1b_3/NOR_0/w_n27_1# ALU_1b_3/NOR_2/A 0.03fF
C82 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# vdd 0.14fF
C83 ALU_1b_3/AND_15/A ALU_1b_3/AND_12/w_64_45# 0.36fF
C84 ALU_1b_2/AND_18/a_78_51# ALU_1b_2/NOR_3/A 0.07fF
C85 ALU_1b_1/AND_4/w_64_45# B3 0.10fF
C86 ALU_1b_2/NOT_6/in gnd 0.07fF
C87 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/full_adder_1/half_adder_1/A 0.14fF
C88 vdd ALU_1b_3/AND_7/w_64_45# 0.14fF
C89 vdd ALU_1b_3/comparator_0/NOR_3/out 0.03fF
C90 C0 ALU_1b_0/AND_8/out 0.01fF
C91 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_3/AND_5/out 0.04fF
C92 ALU_1b_0/NOR_3/B gnd 0.23fF
C93 ALU_1b_0/comparator_0/NOR_0/A ALU_1b_0/comparator_0/NOR_0/out 0.03fF
C94 vdd ALU_1b_2/AND_19/w_64_45# 0.15fF
C95 ALU_1b_2/NOT_1/in ALU_1b_2/AND_5/out 0.21fF
C96 ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.10fF
C97 gnd ALU_1b_3/AND_7/a_78_51# 0.07fF
C98 ALU_1b_3/comparator_0/NOR_0/A ALU_1b_3/comparator_0/NOR_0/B 0.33fF
C99 S1 ALU_1b_2/decoder_0/AND_0/a_78_51# 0.02fF
C100 ALU_1b_0/NOT_1/in ALU_1b_0/NOT_1/w_n36_43# 0.06fF
C101 gnd ALU_1b_2/AND_19/a_78_51# 0.07fF
C102 ALU_1b_0/NOT_5/in ALU_1b_0/NOR_3/B 0.15fF
C103 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/w_n39_45# 0.11fF
C104 ALU_1b_3/decoder_0/AND_2/a_78_51# ALU_1b_3/AND_12/w_64_45# 0.09fF
C105 ALU_1b_1/AND_2/out ALU_1b_1/AND_2/B 0.38fF
C106 ALU_1b_3/AND_6/w_64_45# ALU_1b_3/AND_2/B 0.03fF
C107 ALU_1b_0/AND_3/w_64_45# ALU_1b_0/AND_3/a_78_51# 0.09fF
C108 vdd ALU_1b_3/comparator_0/AND_2/a_78_51# 0.06fF
C109 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.14fF
C110 C1 ALU_1b_0/AND_9/a_78_51# 0.19fF
C111 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_15/B 0.03fF
C112 ALU_1b_0/AND_13/a_78_51# ALU_1b_0/AND_14/B 0.10fF
C113 ALU_1b_1/AND_4/out ALU_1b_1/AND_5/a_78_51# 0.24fF
C114 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C115 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out gnd 0.04fF
C116 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/NOR_0/B 0.01fF
C117 ALU_1b_3/comparator_0/NOR_1/A ALU_1b_3/comparator_0/w_113_n67# 0.06fF
C118 ALU_1b_3/comparator_0/AND_5/a_78_51# ALU_1b_3/AND_7/out 0.14fF
C119 ALU_1b_1/AND_8/out ALU_1b_1/comparator_0/AND_4/a_78_51# 0.20fF
C120 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_14/B 0.06fF
C121 ALU_1b_1/AND_15/B ALU_1b_1/AND_15/A 0.28fF
C122 ALU_1b_3/decoder_0/AND_2/a_78_51# ALU_1b_3/AND_5/B 0.05fF
C123 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.06fF
C124 ALU_1b_1/AND_6/w_64_45# ALU_1b_1/decoder_0/AND_2/B 0.09fF
C125 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C126 vdd ALU_1b_3/comparator_0/AND_4/w_64_45# 0.14fF
C127 ALU_1b_2/AND_1/w_64_45# ALU_1b_2/AND_2/B 0.06fF
C128 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/AND_5/out 0.19fF
C129 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_1/AND_3/out 0.13fF
C130 ALU_1b_2/AND_15/a_78_51# ALU_1b_2/AND_15/A 0.05fF
C131 ALU_1b_3/NOR_4/w_n27_1# ALU_1b_3/NOR_3/A 0.06fF
C132 gnd ALU_1b_3/comparator_0/AND_4/a_78_51# 0.07fF
C133 ALU_1b_0/decoder_0/AND_0/a_78_51# gnd 0.07fF
C134 ALU_1b_2/AND_18/A ALU_1b_2/AND_5/B 0.26fF
C135 vdd ALU_1b_1/comparator_0/w_113_n67# 0.12fF
C136 vdd ALU_1b_2/AND_4/a_78_51# 0.06fF
C137 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_1/A 0.01fF
C138 ALU_1b_1/AND_14/a_78_51# vdd 0.06fF
C139 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.13fF
C140 gnd ALU_1b_3/full_adder_0/half_adder_1/A 0.03fF
C141 ALU_1b_2/comparator_0/w_113_n67# ALU_1b_2/comparator_0/NOR_1/B 0.62fF
C142 ALU_1b_2/full_adder_1/NOR_0/B vdd 0.91fF
C143 ALU_1b_1/AND_0/w_64_45# vdd 0.15fF
C144 ALU_1b_0/NOR_4/A ALU_1b_0/AND_9/w_64_45# 0.03fF
C145 ALU_1b_2/AND_14/a_78_51# ALU_1b_2/AND_15/B 0.05fF
C146 ALU_1b_0/AND_6/out gnd 0.07fF
C147 ALU_1b_2/AND_19/A ALU_1b_2/AND_5/B 0.26fF
C148 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_2/a_n14_7# 0.00fF
C149 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/full_adder_1/half_adder_0/w_36_45# 0.09fF
C150 ALU_1b_3/AND_7/out ALU_1b_3/comparator_0/w_n39_45# 0.06fF
C151 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/AND_1/out 0.06fF
C152 gnd ALU_1b_3/AND_18/A 0.27fF
C153 ALU_1b_1/AND_17/w_64_45# vdd 0.15fF
C154 vdd ALU_1b_1/comparator_0/w_n74_45# 0.06fF
C155 ALU_1b_0/full_adder_1/NOR_0/A ALU_1b_0/full_adder_1/NOR_0/B 0.38fF
C156 ALU_1b_0/NOR_4/B vdd 0.03fF
C157 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.09fF
C158 ALU_1b_2/AND_16/A ALU_1b_2/AND_16/w_64_45# 0.06fF
C159 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_9/out 0.19fF
C160 gnd ALU_1b_2/AND_6/a_78_51# 0.07fF
C161 ALU_1b_0/decoder_0/AND_2/a_78_51# S0 0.05fF
C162 ALU_1b_0/NOR_2/B vdd 0.03fF
C163 ALU_1b_1/AND_17/a_78_51# gnd 0.07fF
C164 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# 0.03fF
C165 ALU_1b_0/comparator_0/NOR_0/A vdd 0.03fF
C166 ALU_1b_3/NOT_6/in ALU_1b_3/NOR_1/A 0.37fF
C167 ALU_1b_1/AND_11/a_78_51# ALU_1b_1/AND_11/B 0.19fF
C168 ALU_1b_0/NOT_6/in gnd 0.07fF
C169 ALU_1b_0/AND_3/w_64_45# ALU_1b_0/AND_3/A 0.09fF
C170 B2 ALU_1b_3/AND_5/B 0.28fF
C171 vdd ALU_1b_3/AND_2/a_78_51# 0.06fF
C172 gnd ALU_1b_3/NOR_4/B 0.07fF
C173 gnd ALU_1b_3/AND_19/A 0.07fF
C174 vdd ALU_1b_2/comparator_0/AND_1/a_78_51# 0.06fF
C175 ALU_1b_2/AND_8/out B1 0.01fF
C176 A0 ALU_1b_0/AND_6/a_78_51# 0.19fF
C177 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.00fF
C178 ALU_1b_1/full_adder_1/half_adder_1/A gnd 0.03fF
C179 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/NOR_0/B 0.38fF
C180 ALU_1b_3/AND_16/w_64_45# ALU_1b_3/AND_16/a_78_51# 0.09fF
C181 ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/AND_11/B 0.05fF
C182 ALU_1b_1/NOR_4/A ALU_1b_1/NOR_4/B 0.35fF
C183 ALU_1b_0/AND_6/w_64_45# ALU_1b_0/decoder_0/AND_1/B 0.13fF
C184 ALU_1b_1/comparator_0/AND_0/w_64_45# ALU_1b_1/comparator_0/NOR_0/A 0.03fF
C185 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_0/a_78_51# 0.29fF
C186 ALU_1b_2/AND_0/w_64_45# ALU_1b_2/AND_0/out 0.09fF
C187 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.06fF
C188 ALU_1b_0/comparator_0/AND_5/B vdd 0.03fF
C189 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/AND_4/out 0.20fF
C190 vdd ALU_1b_3/NOR_0/A 0.20fF
C191 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/half_adder_1/w_36_45# 0.09fF
C192 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_0/NOR_0/B 0.00fF
C193 ALU_1b_2/AND_6/out ALU_1b_2/AND_9/out 0.29fF
C194 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_5/B 0.16fF
C195 ALU_1b_0/AND_9/A ALU_1b_0/AND_6/w_64_45# 0.36fF
C196 ALU_1b_0/comparator_0/NOR_2/A gnd 0.24fF
C197 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/AND_5/out 0.05fF
C198 vdd ALU_1b_2/comparator_0/AND_5/w_64_45# 0.13fF
C199 ALU_1b_0/AND_9/w_64_45# C1 0.06fF
C200 ALU_1b_2/NOR_1/B ALU_1b_2/C0 0.01fF
C201 ALU_1b_0/AND_16/w_64_45# ALU_1b_0/AND_2/B 0.10fF
C202 ALU_1b_1/AND_19/w_64_45# ALU_1b_1/AND_19/A 0.06fF
C203 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out 0.09fF
C204 Cout gnd 0.07fF
C205 vdd ALU_1b_3/AND_2/out 0.35fF
C206 ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/AND_2/w_64_45# 0.16fF
C207 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_5/w_64_45# 0.03fF
C208 gnd ALU_1b_2/comparator_0/AND_5/a_78_51# 0.07fF
C209 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.01fF
C210 ALU_1b_1/AND_5/a_78_51# vdd 0.06fF
C211 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/NOR_1/A 0.03fF
C212 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/NOR_0/B 0.48fF
C213 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_0/AND_4/out 0.06fF
C214 ALU_1b_0/AND_9/a_78_51# vdd 0.06fF
C215 ALU_1b_1/NOR_2/A ALU_1b_1/NOT_3/in 0.23fF
C216 ALU_1b_0/AND_17/A ALU_1b_0/AND_17/a_78_51# 0.03fF
C217 ALU_1b_3/AND_0/out ALU_1b_3/AND_2/a_78_51# 0.10fF
C218 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_1/A 0.11fF
C219 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out gnd 0.04fF
C220 ALU_1b_0/NOR_0/B ALU_1b_0/NOR_3/A 0.01fF
C221 ALU_1b_0/comparator_0/NOR_0/B gnd 0.17fF
C222 ALU_1b_1/AND_0/out B3 0.01fF
C223 vdd ALU_1b_2/AND_14/A 0.03fF
C224 S1 ALU_1b_3/AND_12/w_64_45# 0.06fF
C225 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/AND_5/out 0.02fF
C226 ALU_1b_1/AND_19/a_78_51# ALU_1b_1/NOR_0/A 0.16fF
C227 ALU_1b_3/AND_2/out ALU_1b_3/AND_1/a_78_51# 0.24fF
C228 vdd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.22fF
C229 Cin ALU_1b_0/AND_2/B 0.27fF
C230 vdd ALU_1b_1/decoder_0/AND_2/B 0.03fF
C231 ALU_1b_0/AND_5/out ALU_1b_0/AND_5/w_64_45# 0.03fF
C232 ALU_1b_0/AND_16/w_64_45# vdd 0.15fF
C233 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.13fF
C234 ALU_1b_0/AND_4/out C0 0.01fF
C235 ALU_1b_1/AND_11/a_78_51# gnd 0.07fF
C236 ALU_1b_2/AND_7/w_64_45# ALU_1b_2/AND_7/out 0.03fF
C237 vdd ALU_1b_3/comparator_0/NOR_2/B 0.31fF
C238 ALU_1b_0/full_adder_0/w_448_45# ALU_1b_0/full_adder_0/NOR_0/B 0.16fF
C239 ALU_1b_1/AND_11/B gnd 0.13fF
C240 ALU_1b_1/AND_12/w_64_45# ALU_1b_1/AND_5/B 0.03fF
C241 ALU_1b_2/AND_5/out ALU_1b_2/C0 0.01fF
C242 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.05fF
C243 ALU_1b_0/AND_16/a_78_51# gnd 0.07fF
C244 ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.26fF
C245 vdd ALU_1b_2/comparator_0/NOR_1/out 0.03fF
C246 S1 ALU_1b_3/AND_5/B 0.03fF
C247 ALU_1b_0/AND_9/A ALU_1b_0/AND_10/B 0.29fF
C248 ALU_1b_3/AND_2/out ALU_1b_3/AND_0/out 0.96fF
C249 gnd ALU_1b_3/comparator_0/NOR_2/out 0.07fF
C250 ALU_1b_1/comparator_0/AND_0/a_78_51# vdd 0.06fF
C251 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.03fF
C252 ALU_1b_3/AND_8/w_64_45# ALU_1b_3/AND_8/a_78_51# 0.09fF
C253 ALU_1b_3/AND_11/a_78_51# ALU_1b_3/AND_9/A 0.03fF
C254 ALU_1b_3/AND_9/A ALU_1b_3/AND_11/B 0.37fF
C255 ALU_1b_1/AND_3/a_78_51# ALU_1b_1/AND_3/A 0.03fF
C256 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.06fF
C257 ALU_1b_2/AND_4/out ALU_1b_2/full_adder_1/half_adder_1/A 0.11fF
C258 vdd ALU_1b_3/NOT_1/w_n36_43# 0.06fF
C259 ALU_1b_1/NOR_2/A ALU_1b_1/NOR_2/w_n27_1# 0.06fF
C260 ALU_1b_0/comparator_0/AND_3/a_78_51# ALU_1b_0/AND_8/out 0.03fF
C261 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_4/a_78_51# 0.04fF
C262 Cin vdd 0.19fF
C263 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.00fF
C264 ALU_1b_3/AND_12/w_64_45# ALU_1b_3/decoder_0/AND_1/B 0.03fF
C265 vdd ALU_1b_2/NOR_3/B 0.33fF
C266 ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C267 ALU_1b_2/AND_14/B ALU_1b_2/AND_12/w_64_45# 0.03fF
C268 ALU_1b_3/comparator_0/AND_3/w_64_45# ALU_1b_3/AND_8/out 0.16fF
C269 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out gnd 0.04fF
C270 ALU_1b_2/AND_4/a_78_51# B1 0.03fF
C271 S0 ALU_1b_2/decoder_0/AND_2/B 0.29fF
C272 ALU_1b_0/decoder_0/AND_1/a_78_51# ALU_1b_0/decoder_0/AND_1/B 0.19fF
C273 ALU_1b_1/comparator_0/AND_3/w_64_45# vdd 0.15fF
C274 ALU_1b_3/NOT_6/in ALU_1b_3/NOR_4/w_n27_1# 0.11fF
C275 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_14/A 0.09fF
C276 ALU_1b_2/NOR_4/w_n27_1# ALU_1b_2/NOR_3/B 0.20fF
C277 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_74# vdd 0.02fF
C278 ALU_1b_1/AND_2/w_64_45# vdd 0.15fF
C279 ALU_1b_1/comparator_0/AND_3/a_78_51# gnd 0.07fF
C280 ALU_1b_2/comparator_0/AND_4/w_64_45# ALU_1b_2/AND_7/out 0.10fF
C281 ALU_1b_1/AND_4/out ALU_1b_1/C0 0.16fF
C282 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_0/half_adder_1/A 0.26fF
C283 ALU_1b_2/AND_14/A ALU_1b_2/AND_15/A 0.10fF
C284 ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/AND_2/B 0.05fF
C285 ALU_1b_3/full_adder_1/NOR_0/out ALU_1b_3/AND_18/A 0.04fF
C286 ALU_1b_0/decoder_0/AND_1/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C287 ALU_1b_1/AND_5/B gnd 0.48fF
C288 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_0/full_adder_0/NOR_0/B 0.00fF
C289 vdd ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out 0.06fF
C290 ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/w_n39_45# 0.15fF
C291 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# vdd 0.22fF
C292 vdd ALU_1b_1/NOR_2/w_n27_1# 0.24fF
C293 gnd ALU_1b_3/full_adder_0/NOR_0/B 0.07fF
C294 ALU_1b_0/AND_9/w_64_45# vdd 0.42fF
C295 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/w_n74_45# 0.03fF
C296 ALU_1b_2/AND_8/out ALU_1b_2/AND_9/A 0.12fF
C297 ALU_1b_0/AND_3/out ALU_1b_0/AND_5/a_78_51# 0.10fF
C298 C1 ALU_1b_0/NOR_1/B 0.01fF
C299 ALU_1b_0/AND_19/w_64_45# ALU_1b_0/AND_5/B 0.06fF
C300 ALU_1b_0/AND_10/a_78_51# gnd 0.07fF
C301 gnd ALU_1b_3/AND_14/B 0.07fF
C302 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.06fF
C303 vdd ALU_1b_2/decoder_0/AND_0/a_78_51# 0.06fF
C304 ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/NOR_0/out 0.15fF
C305 ALU_1b_1/AND_7/out ALU_1b_1/comparator_0/w_n74_45# 0.10fF
C306 ALU_1b_3/AND_14/A ALU_1b_3/AND_14/a_78_51# 0.03fF
C307 ALU_1b_1/AND_15/B ALU_1b_1/AND_15/w_64_45# 0.06fF
C308 ALU_1b_2/AND_0/out ALU_1b_2/AND_2/w_64_45# 0.20fF
C309 ALU_1b_1/NOR_1/B ALU_1b_1/NOR_1/A 0.33fF
C310 ALU_1b_0/NOT_5/in gnd 0.07fF
C311 ALU_1b_1/comparator_0/w_n220_n67# ALU_1b_1/comparator_0/NOR_2/B 0.62fF
C312 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_10/a_78_51# 0.09fF
C313 ALU_1b_3/AND_3/a_78_51# ALU_1b_3/AND_5/B 0.29fF
C314 ALU_1b_3/NOT_1/in ALU_1b_3/NOT_1/w_n36_43# 0.06fF
C315 ALU_1b_2/AND_3/out gnd 0.11fF
C316 ALU_1b_0/comparator_0/NOR_3/B vdd 0.03fF
C317 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/NOR_0/B 0.00fF
C318 ALU_1b_2/AND_15/w_64_45# ALU_1b_2/AND_15/a_78_51# 0.09fF
C319 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_2/AND_5/out 0.10fF
C320 ALU_1b_0/decoder_0/AND_1/B S0 0.03fF
C321 ALU_1b_3/AND_16/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.03fF
C322 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/NOR_3/B 0.43fF
C323 ALU_1b_0/comparator_0/NOR_3/out gnd 0.07fF
C324 vdd ALU_1b_2/AND_6/out 0.20fF
C325 ALU_1b_3/comparator_0/w_113_n67# ALU_1b_3/comparator_0/NOR_1/out 0.11fF
C326 ALU_1b_0/AND_7/out B0 0.28fF
C327 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/w_448_45# 0.06fF
C328 ALU_1b_1/NOR_0/B vdd 0.20fF
C329 ALU_1b_3/full_adder_0/half_adder_1/w_36_45# ALU_1b_3/full_adder_0/half_adder_1/A 0.06fF
C330 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# vdd 0.14fF
C331 gnd ALU_1b_2/decoder_0/AND_3/a_78_51# 0.07fF
C332 ALU_1b_0/comparator_0/AND_2/w_64_45# vdd 0.15fF
C333 ALU_1b_1/AND_1/out vdd 0.35fF
C334 vdd ALU_1b_3/AND_17/a_78_51# 0.06fF
C335 ALU_1b_1/AND_1/w_64_45# ALU_1b_1/AND_1/a_78_51# 0.09fF
C336 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/full_adder_0/NOR_0/B 0.15fF
C337 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/NOR_0/B 0.48fF
C338 ALU_1b_2/comparator_0/AND_0/w_64_45# ALU_1b_2/AND_6/out 0.26fF
C339 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_2/AND_16/A 0.03fF
C340 ALU_1b_3/AND_16/A ALU_1b_3/AND_16/a_78_51# 0.03fF
C341 ALU_1b_0/comparator_0/AND_0/w_64_45# ALU_1b_0/AND_9/out 0.30fF
C342 ALU_1b_0/comparator_0/AND_2/a_78_51# gnd 0.07fF
C343 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.09fF
C344 vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.02fF
C345 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/AND_5/out 0.02fF
C346 ALU_1b_0/AND_4/a_78_51# ALU_1b_0/AND_5/B 0.29fF
C347 ALU_1b_1/AND_8/out ALU_1b_1/AND_6/w_64_45# 0.15fF
C348 ALU_1b_2/AND_4/out ALU_1b_2/AND_5/B 0.38fF
C349 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/NOR_3/out 0.15fF
C350 ALU_1b_1/AND_1/w_64_45# ALU_1b_1/AND_0/out 0.20fF
C351 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd 0.06fF
C352 ALU_1b_1/NOR_3/A gnd 0.23fF
C353 vdd ALU_1b_3/full_adder_0/NOR_0/A 0.03fF
C354 ALU_1b_3/AND_4/w_64_45# ALU_1b_3/AND_5/B 0.06fF
C355 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/NOR_0/B 0.09fF
C356 ALU_1b_2/AND_1/out ALU_1b_2/AND_1/a_78_51# 0.05fF
C357 ALU_1b_2/NOT_3/in ALU_1b_2/NOR_2/B 0.03fF
C358 ALU_1b_0/AND_17/a_78_51# ALU_1b_0/NOR_3/B 0.07fF
C359 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/AND_4/out 0.09fF
C360 ALU_1b_2/comparator_0/AND_0/a_78_51# ALU_1b_2/comparator_0/NOR_0/A 0.05fF
C361 ALU_1b_2/NOT_6/in ALU_1b_2/NOR_4/B 0.15fF
C362 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_2/A 0.33fF
C363 vdd ALU_1b_2/comparator_0/NOR_2/A 0.03fF
C364 ALU_1b_3/AND_17/w_64_45# ALU_1b_3/NOR_3/B 0.07fF
C365 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/w_36_45# 0.03fF
C366 vdd ALU_1b_1/C0 0.56fF
C367 gnd F0 0.50fF
C368 ALU_1b_1/NOT_4/in ALU_1b_1/NOR_2/w_n27_1# 0.11fF
C369 gnd ALU_1b_3/AND_4/out 0.07fF
C370 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C371 ALU_1b_2/AND_1/out ALU_1b_2/AND_0/out 0.11fF
C372 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_2/full_adder_1/half_adder_1/A 0.03fF
C373 ALU_1b_3/AND_3/A ALU_1b_3/AND_5/B 0.42fF
C374 ALU_1b_1/AND_16/a_78_51# ALU_1b_1/AND_2/B 0.19fF
C375 ALU_1b_2/AND_3/out ALU_1b_2/AND_3/w_64_45# 0.09fF
C376 ALU_1b_2/AND_19/A ALU_1b_2/AND_19/a_78_51# 0.03fF
C377 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/NOT_1/in 0.06fF
C378 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C379 ALU_1b_2/AND_17/A gnd 0.34fF
C380 ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/AND_2/a_78_51# 0.03fF
C381 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_5/a_78_51# 0.05fF
C382 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_4/a_78_51# 0.18fF
C383 ALU_1b_0/NOT_2/in ALU_1b_0/NOR_0/w_n27_1# 0.11fF
C384 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C385 ALU_1b_2/AND_10/a_78_51# ALU_1b_2/NOR_1/A 0.05fF
C386 vdd ALU_1b_2/comparator_0/NOR_0/B 0.09fF
C387 vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.02fF
C388 ALU_1b_2/AND_3/out F0 0.01fF
C389 ALU_1b_1/AND_18/w_64_45# ALU_1b_1/AND_18/a_78_51# 0.09fF
C390 ALU_1b_2/AND_12/a_78_51# ALU_1b_2/AND_12/w_64_45# 0.09fF
C391 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/AND_7/out 0.11fF
C392 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_4/w_64_45# 0.03fF
C393 ALU_1b_3/comparator_0/AND_2/w_64_45# ALU_1b_3/comparator_0/AND_2/a_78_51# 0.09fF
C394 ALU_1b_1/NOT_6/in Cout 0.03fF
C395 ALU_1b_1/comparator_0/w_n195_n67# vdd 0.12fF
C396 gnd ALU_1b_2/comparator_0/NOR_0/out 0.07fF
C397 ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.26fF
C398 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C399 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C400 ALU_1b_0/NOR_1/B vdd 0.20fF
C401 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/NOR_0/out 0.03fF
C402 ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C403 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C404 ALU_1b_2/comparator_0/AND_3/w_64_45# ALU_1b_2/comparator_0/AND_5/B 0.06fF
C405 ALU_1b_2/NOR_2/B ALU_1b_2/NOR_2/w_n27_1# 0.09fF
C406 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_3/NOT_1/in 0.03fF
C407 vdd ALU_1b_3/AND_11/a_78_51# 0.06fF
C408 vdd ALU_1b_3/AND_11/B 1.14fF
C409 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_2/AND_5/out 0.04fF
C410 ALU_1b_0/AND_2/a_78_51# gnd 0.07fF
C411 ALU_1b_0/AND_4/out ALU_1b_0/AND_5/B 0.38fF
C412 vdd ALU_1b_2/AND_16/a_78_51# 0.06fF
C413 ALU_1b_3/AND_2/out ALU_1b_3/C0 0.16fF
C414 ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/AND_10/B 0.09fF
C415 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/NOR_0/out 0.15fF
C416 ALU_1b_3/NOT_1/in ALU_1b_3/full_adder_1/half_adder_1/A 0.23fF
C417 gnd ALU_1b_3/comparator_0/AND_2/B 0.07fF
C418 ALU_1b_2/AND_5/a_78_51# ALU_1b_2/C0 0.03fF
C419 ALU_1b_1/AND_5/out ALU_1b_1/AND_5/w_64_45# 0.03fF
C420 ALU_1b_3/AND_7/a_78_51# ALU_1b_3/AND_7/out 0.16fF
C421 gnd ALU_1b_3/AND_10/B 0.13fF
C422 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_4/a_78_8# 0.00fF
C423 ALU_1b_2/full_adder_1/w_448_45# vdd 0.12fF
C424 ALU_1b_0/AND_0/out C1 0.01fF
C425 F3 ALU_1b_1/NOR_2/w_n27_1# 0.03fF
C426 gnd ALU_1b_3/full_adder_1/NOR_0/out 0.07fF
C427 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_0/NOR_0/B 0.00fF
C428 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C429 ALU_1b_2/AND_0/a_78_51# gnd 0.07fF
C430 ALU_1b_0/decoder_0/AND_2/B S1 0.07fF
C431 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/w_36_45# 0.12fF
C432 ALU_1b_0/NOR_0/A gnd 0.17fF
C433 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/w_36_45# 0.29fF
C434 vdd ALU_1b_2/AND_18/w_64_45# 0.15fF
C435 vdd ALU_1b_3/AND_12/w_64_45# 0.47fF
C436 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_2/C0 0.03fF
C437 ALU_1b_0/full_adder_1/NOR_0/A vdd 0.03fF
C438 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C439 gnd ALU_1b_3/AND_12/a_78_51# 0.07fF
C440 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.20fF
C441 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/w_n74_45# 0.18fF
C442 gnd ALU_1b_2/AND_18/a_78_51# 0.07fF
C443 vdd ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.06fF
C444 ALU_1b_1/AND_3/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.26fF
C445 ALU_1b_1/comparator_0/NOR_1/A vdd 0.03fF
C446 ALU_1b_3/AND_12/a_78_51# ALU_1b_3/AND_14/B 0.05fF
C447 gnd ALU_1b_3/NOR_2/A 0.07fF
C448 gnd ALU_1b_2/AND_2/B 0.48fF
C449 vdd ALU_1b_3/comparator_0/AND_3/a_78_51# 0.06fF
C450 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out 0.05fF
C451 ALU_1b_2/comparator_0/NOR_1/A ALU_1b_2/comparator_0/NOR_1/B 0.33fF
C452 ALU_1b_0/AND_7/out ALU_1b_0/AND_9/A 0.01fF
C453 ALU_1b_2/NOR_4/A ALU_1b_2/AND_9/w_64_45# 0.03fF
C454 ALU_1b_2/AND_13/a_78_51# ALU_1b_2/AND_14/A 0.05fF
C455 ALU_1b_1/AND_4/out ALU_1b_1/AND_4/a_78_51# 0.05fF
C456 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.09fF
C457 vdd ALU_1b_3/AND_5/B 0.10fF
C458 ALU_1b_2/AND_4/w_64_45# ALU_1b_2/AND_4/a_78_51# 0.09fF
C459 gnd ALU_1b_3/decoder_0/AND_1/a_78_51# 0.07fF
C460 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.52fF
C461 ALU_1b_3/AND_7/out ALU_1b_3/comparator_0/AND_4/a_78_51# 0.03fF
C462 ALU_1b_0/AND_1/out gnd 0.69fF
C463 ALU_1b_1/AND_8/out vdd 0.66fF
C464 A0 ALU_1b_0/AND_2/B 0.50fF
C465 ALU_1b_1/AND_14/A ALU_1b_1/AND_14/B 0.42fF
C466 ALU_1b_1/AND_9/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C467 ALU_1b_1/full_adder_1/NOR_0/B vdd 0.91fF
C468 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_74# 0.01fF
C469 ALU_1b_3/AND_3/out ALU_1b_3/AND_5/w_64_45# 0.20fF
C470 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.09fF
C471 vdd ALU_1b_3/comparator_0/w_88_n67# 0.12fF
C472 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# ALU_1b_1/full_adder_0/NOR_0/B 0.12fF
C473 ALU_1b_0/AND_0/a_78_51# ALU_1b_0/AND_2/B 0.14fF
C474 ALU_1b_0/comparator_0/NOR_2/B gnd 0.07fF
C475 ALU_1b_3/comparator_0/w_88_n67# ALU_1b_3/comparator_0/NOR_1/B 0.19fF
C476 ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/w_113_n67# 0.02fF
C477 vdd ALU_1b_2/AND_10/a_78_51# 0.06fF
C478 ALU_1b_1/AND_15/a_78_51# vdd 0.06fF
C479 ALU_1b_1/NOR_0/A ALU_1b_1/NOR_0/w_n27_1# 0.06fF
C480 ALU_1b_3/full_adder_0/half_adder_1/w_36_45# ALU_1b_3/full_adder_0/NOR_0/B 0.36fF
C481 ALU_1b_1/NOR_4/A vdd 0.10fF
C482 gnd ALU_1b_2/comparator_0/NOR_3/A 0.21fF
C483 ALU_1b_1/full_adder_0/NOR_0/A gnd 0.07fF
C484 ALU_1b_1/AND_19/a_78_51# ALU_1b_1/AND_5/B 0.19fF
C485 ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/decoder_0/AND_2/B 0.03fF
C486 A0 vdd 0.21fF
C487 ALU_1b_1/comparator_0/w_n220_n67# ALU_1b_1/AND_11/B 0.03fF
C488 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C489 ALU_1b_0/AND_0/out ALU_1b_0/AND_2/B 0.11fF
C490 ALU_1b_2/AND_15/B ALU_1b_2/AND_15/a_78_51# 0.19fF
C491 ALU_1b_2/comparator_0/w_n220_n67# ALU_1b_2/comparator_0/NOR_2/out 0.11fF
C492 ALU_1b_1/NOT_6/in gnd 0.07fF
C493 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_3/out 0.05fF
C494 vdd ALU_1b_2/AND_7/w_64_45# 0.14fF
C495 vdd ALU_1b_2/comparator_0/NOR_3/out 0.03fF
C496 ALU_1b_1/AND_19/w_64_45# vdd 0.15fF
C497 ALU_1b_0/AND_0/a_78_51# vdd 0.06fF
C498 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C499 ALU_1b_0/AND_2/w_64_45# ALU_1b_0/AND_2/a_78_51# 0.09fF
C500 gnd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# 0.02fF
C501 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.01fF
C502 gnd ALU_1b_2/AND_7/a_78_51# 0.07fF
C503 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/NOR_3/out 0.03fF
C504 S1 ALU_1b_1/decoder_0/AND_0/a_78_51# 0.02fF
C505 ALU_1b_1/AND_19/a_78_51# gnd 0.07fF
C506 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.01fF
C507 ALU_1b_1/full_adder_1/w_448_45# ALU_1b_1/AND_18/A 0.03fF
C508 ALU_1b_2/AND_16/w_64_45# ALU_1b_2/NOR_0/B 0.03fF
C509 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# 0.03fF
C510 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/AND_5/out 0.06fF
C511 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C512 C0 gnd 0.31fF
C513 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/NOR_0/A 0.12fF
C514 vdd ALU_1b_2/comparator_0/AND_2/a_78_51# 0.06fF
C515 ALU_1b_0/AND_0/out vdd 0.03fF
C516 F0 ALU_1b_2/AND_2/B 0.01fF
C517 ALU_1b_1/AND_0/out ALU_1b_1/AND_1/a_78_51# 0.10fF
C518 ALU_1b_1/AND_18/A ALU_1b_1/AND_18/w_64_45# 0.06fF
C519 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/AND_4/out 0.06fF
C520 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_0/a_78_51# 0.14fF
C521 ALU_1b_3/decoder_0/AND_1/a_78_51# ALU_1b_3/AND_6/w_64_45# 0.09fF
C522 ALU_1b_1/comparator_0/AND_0/a_78_51# ALU_1b_1/AND_9/out 0.02fF
C523 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_1/a_78_51# 0.10fF
C524 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C525 ALU_1b_1/AND_7/w_64_45# ALU_1b_1/AND_7/a_78_51# 0.09fF
C526 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# ALU_1b_1/full_adder_1/NOR_0/A 0.03fF
C527 ALU_1b_2/AND_17/A ALU_1b_2/AND_2/B 0.26fF
C528 ALU_1b_1/NOR_1/B B3 0.01fF
C529 vdd ALU_1b_3/NOR_3/A 0.22fF
C530 ALU_1b_0/AND_19/w_64_45# ALU_1b_0/AND_19/a_78_51# 0.09fF
C531 ALU_1b_2/comparator_0/AND_1/w_64_45# ALU_1b_2/comparator_0/AND_1/a_78_51# 0.09fF
C532 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C533 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C534 vdd ALU_1b_2/comparator_0/AND_4/w_64_45# 0.14fF
C535 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/AND_3/out 0.14fF
C536 ALU_1b_0/AND_17/w_64_45# ALU_1b_0/AND_2/B 0.06fF
C537 ALU_1b_0/NOR_2/A ALU_1b_0/NOR_2/B 0.47fF
C538 ALU_1b_1/AND_2/out vdd 0.35fF
C539 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.26fF
C540 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_3/AND_16/A 0.03fF
C541 ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/decoder_0/AND_1/B 0.29fF
C542 gnd ALU_1b_2/comparator_0/AND_4/a_78_51# 0.07fF
C543 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/w_448_45# 0.06fF
C544 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOR_1/A 0.09fF
C545 ALU_1b_0/comparator_0/w_113_n67# vdd 0.12fF
C546 ALU_1b_1/AND_4/a_78_51# vdd 0.06fF
C547 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_9/A 0.95fF
C548 A3 ALU_1b_1/AND_15/A 0.42fF
C549 ALU_1b_2/AND_1/out ALU_1b_2/C0 0.01fF
C550 ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/comparator_0/NOR_2/A 0.03fF
C551 ALU_1b_0/AND_14/a_78_51# vdd 0.06fF
C552 ALU_1b_1/AND_2/a_78_51# ALU_1b_1/AND_2/B 0.29fF
C553 ALU_1b_0/NOR_3/B ALU_1b_0/NOR_3/A 0.34fF
C554 ALU_1b_2/full_adder_0/half_adder_1/A gnd 0.03fF
C555 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_8/out 0.11fF
C556 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.06fF
C557 vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.06fF
C558 gnd ALU_1b_3/NOT_4/in 0.07fF
C559 ALU_1b_0/full_adder_0/NOR_0/B vdd 0.91fF
C560 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.03fF
C561 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.01fF
C562 ALU_1b_1/NOR_1/A ALU_1b_1/NOT_3/in 0.03fF
C563 ALU_1b_3/decoder_0/AND_3/a_78_51# ALU_1b_3/AND_15/A 0.05fF
C564 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_4/B 0.03fF
C565 ALU_1b_3/AND_1/w_64_45# vdd 0.15fF
C566 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_4/a_78_8# 0.00fF
C567 gnd ALU_1b_2/AND_18/A 0.27fF
C568 ALU_1b_0/AND_17/w_64_45# vdd 0.15fF
C569 ALU_1b_0/comparator_0/w_n74_45# vdd 0.06fF
C570 ALU_1b_2/AND_0/a_78_51# ALU_1b_2/AND_2/B 0.14fF
C571 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out 0.08fF
C572 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# vdd 0.14fF
C573 ALU_1b_1/AND_6/a_78_51# gnd 0.07fF
C574 ALU_1b_2/AND_6/out ALU_1b_2/AND_9/A 0.01fF
C575 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_3/AND_5/out 0.05fF
C576 ALU_1b_0/AND_8/w_64_45# ALU_1b_0/AND_8/out 0.03fF
C577 ALU_1b_0/AND_17/a_78_51# gnd 0.07fF
C578 ALU_1b_0/comparator_0/AND_3/a_78_51# ALU_1b_0/comparator_0/NOR_2/A 0.17fF
C579 ALU_1b_0/AND_9/out ALU_1b_0/AND_9/A 0.04fF
C580 ALU_1b_1/AND_5/B F2 0.01fF
C581 vdd ALU_1b_2/AND_2/a_78_51# 0.06fF
C582 ALU_1b_2/NOR_4/B gnd 0.07fF
C583 ALU_1b_3/comparator_0/NOR_0/A ALU_1b_3/comparator_0/w_88_n67# 0.06fF
C584 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_3/a_78_51# 0.19fF
C585 ALU_1b_3/comparator_0/AND_3/w_64_45# ALU_1b_3/comparator_0/NOR_2/A 0.03fF
C586 ALU_1b_1/comparator_0/AND_1/a_78_51# vdd 0.06fF
C587 ALU_1b_2/AND_0/w_64_45# A1 0.10fF
C588 gnd ALU_1b_2/AND_19/A 0.07fF
C589 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_0/NOR_0/A 0.06fF
C590 ALU_1b_3/AND_1/w_64_45# ALU_1b_3/AND_1/a_78_51# 0.09fF
C591 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C592 ALU_1b_3/full_adder_1/half_adder_1/w_36_45# ALU_1b_3/full_adder_1/NOR_0/B 0.36fF
C593 ALU_1b_1/comparator_0/NOR_1/out ALU_1b_1/AND_10/B 0.05fF
C594 ALU_1b_1/AND_5/w_64_45# ALU_1b_1/AND_5/a_78_51# 0.09fF
C595 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/AND_8/out 0.38fF
C596 ALU_1b_2/NOR_1/B ALU_1b_2/NOT_3/in 0.15fF
C597 ALU_1b_0/comparator_0/AND_5/a_78_51# ALU_1b_0/AND_8/out 0.02fF
C598 vdd ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.06fF
C599 ALU_1b_2/AND_5/out ALU_1b_2/AND_5/a_78_51# 0.05fF
C600 ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C601 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_14/a_78_51# 0.09fF
C602 ALU_1b_0/AND_8/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C603 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_1/AND_4/out 0.70fF
C604 vdd ALU_1b_2/NOR_0/A 0.20fF
C605 ALU_1b_0/full_adder_0/w_448_45# ALU_1b_0/AND_17/A 0.03fF
C606 ALU_1b_1/AND_3/out ALU_1b_1/full_adder_1/half_adder_1/A 0.23fF
C607 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/NOR_0/B 0.48fF
C608 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.05fF
C609 gnd F2 0.50fF
C610 ALU_1b_3/comparator_0/AND_5/w_64_45# ALU_1b_3/AND_8/out 0.32fF
C611 vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.06fF
C612 ALU_1b_3/AND_1/w_64_45# ALU_1b_3/AND_0/out 0.20fF
C613 ALU_1b_1/comparator_0/AND_5/w_64_45# vdd 0.13fF
C614 ALU_1b_1/comparator_0/AND_4/w_64_45# ALU_1b_1/comparator_0/AND_4/a_78_51# 0.09fF
C615 ALU_1b_1/AND_7/out ALU_1b_1/AND_8/out 0.40fF
C616 ALU_1b_3/AND_8/w_64_45# ALU_1b_3/AND_9/A 0.39fF
C617 ALU_1b_1/AND_14/a_78_51# ALU_1b_1/AND_15/A 0.00fF
C618 ALU_1b_1/NOR_1/A ALU_1b_1/NOR_2/w_n27_1# 0.10fF
C619 ALU_1b_2/AND_2/out vdd 0.35fF
C620 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.06fF
C621 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.09fF
C622 ALU_1b_1/AND_6/w_64_45# ALU_1b_1/decoder_0/AND_0/a_78_51# 0.09fF
C623 ALU_1b_1/comparator_0/AND_5/a_78_51# gnd 0.07fF
C624 A3 B3 0.64fF
C625 ALU_1b_3/AND_3/out B2 0.01fF
C626 ALU_1b_0/AND_5/a_78_51# vdd 0.06fF
C627 ALU_1b_0/comparator_0/w_88_n67# ALU_1b_0/comparator_0/NOR_0/B 0.20fF
C628 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/NOT_1/in 0.06fF
C629 ALU_1b_0/NOR_0/B ALU_1b_0/NOR_0/w_n27_1# 0.06fF
C630 ALU_1b_0/NOR_1/A ALU_1b_0/AND_9/A 0.03fF
C631 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# 0.06fF
C632 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out gnd 0.04fF
C633 gnd ALU_1b_3/AND_7/out 0.07fF
C634 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_2/AND_5/out 0.00fF
C635 ALU_1b_2/AND_7/w_64_45# B1 0.06fF
C636 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/NOR_0/B 0.06fF
C637 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# 0.04fF
C638 ALU_1b_3/comparator_0/NOR_1/A ALU_1b_3/comparator_0/NOR_1/out 0.03fF
C639 ALU_1b_1/AND_14/A vdd 0.03fF
C640 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/NOR_0/B 0.00fF
C641 S1 ALU_1b_2/AND_12/w_64_45# 0.06fF
C642 ALU_1b_1/AND_6/out ALU_1b_1/AND_6/w_64_45# 0.14fF
C643 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_0/out 0.23fF
C644 ALU_1b_2/NOT_4/in F1 0.03fF
C645 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# vdd 0.22fF
C646 ALU_1b_0/decoder_0/AND_2/B vdd 0.03fF
C647 ALU_1b_0/AND_3/out ALU_1b_0/AND_4/a_78_51# 0.10fF
C648 ALU_1b_2/NOR_1/B ALU_1b_2/NOR_2/w_n27_1# 0.06fF
C649 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_1/half_adder_1/A 0.26fF
C650 ALU_1b_0/AND_18/w_64_45# ALU_1b_0/AND_5/B 0.10fF
C651 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_6/w_64_45# 0.09fF
C652 ALU_1b_0/AND_11/a_78_51# gnd 0.07fF
C653 ALU_1b_0/AND_11/B gnd 0.13fF
C654 vdd ALU_1b_2/comparator_0/NOR_2/B 0.31fF
C655 ALU_1b_0/AND_15/A B0 0.28fF
C656 vdd ALU_1b_1/comparator_0/NOR_1/out 0.03fF
C657 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_10/B 0.20fF
C658 ALU_1b_3/NOR_0/A ALU_1b_3/NOT_2/in 0.03fF
C659 ALU_1b_1/AND_15/w_64_45# ALU_1b_1/NOR_1/B 0.06fF
C660 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# vdd 0.14fF
C661 S1 ALU_1b_2/AND_5/B 0.03fF
C662 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_11/a_78_51# 0.09fF
C663 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/NOR_0/B 0.38fF
C664 gnd ALU_1b_2/comparator_0/NOR_2/out 0.07fF
C665 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_11/B 0.11fF
C666 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# ALU_1b_0/AND_4/out 0.29fF
C667 ALU_1b_0/comparator_0/AND_0/a_78_51# vdd 0.06fF
C668 ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/comparator_0/NOR_1/out 0.25fF
C669 ALU_1b_1/AND_17/A ALU_1b_1/AND_17/a_78_51# 0.03fF
C670 ALU_1b_3/C0 ALU_1b_3/AND_5/B 0.28fF
C671 ALU_1b_0/NOT_4/in ALU_1b_0/NOR_2/B 0.15fF
C672 ALU_1b_2/comparator_0/w_n195_n67# ALU_1b_2/comparator_0/NOR_3/B 0.06fF
C673 ALU_1b_3/NOR_4/B ALU_1b_3/NOR_1/A 0.07fF
C674 ALU_1b_2/AND_8/out ALU_1b_2/C0 0.01fF
C675 vdd ALU_1b_2/NOT_1/w_n36_43# 0.06fF
C676 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C677 ALU_1b_0/AND_1/out C0 0.01fF
C678 ALU_1b_1/NOR_3/B vdd 0.33fF
C679 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/A 0.16fF
C680 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/C0 0.19fF
C681 ALU_1b_1/comparator_0/AND_0/w_64_45# ALU_1b_1/comparator_0/AND_0/a_78_51# 0.09fF
C682 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_2/B 0.40fF
C683 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_74# 0.01fF
C684 ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.13fF
C685 ALU_1b_1/decoder_0/AND_2/B S0 0.29fF
C686 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/AND_5/out 0.08fF
C687 ALU_1b_0/comparator_0/AND_3/w_64_45# vdd 0.15fF
C688 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/full_adder_1/NOR_0/B 0.15fF
C689 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_74# vdd 0.02fF
C690 vdd ALU_1b_3/AND_19/a_78_51# 0.06fF
C691 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/NOR_0/B 0.01fF
C692 ALU_1b_0/AND_3/w_64_45# A0 0.10fF
C693 ALU_1b_2/AND_1/out ALU_1b_2/AND_16/A 0.11fF
C694 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_1/w_64_45# 0.10fF
C695 ALU_1b_0/comparator_0/AND_1/w_64_45# ALU_1b_0/AND_9/out 0.39fF
C696 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_2/w_64_45# 0.06fF
C697 ALU_1b_0/comparator_0/AND_3/a_78_51# gnd 0.07fF
C698 ALU_1b_1/full_adder_0/w_448_45# ALU_1b_1/full_adder_0/NOR_0/out 0.11fF
C699 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.04fF
C700 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# ALU_1b_0/full_adder_0/half_adder_1/A 0.06fF
C701 ALU_1b_0/AND_5/B gnd 0.48fF
C702 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.03fF
C703 ALU_1b_3/AND_16/a_78_51# ALU_1b_3/NOR_0/B 0.05fF
C704 ALU_1b_3/full_adder_0/half_adder_0/w_36_45# ALU_1b_3/full_adder_0/NOR_0/B 0.12fF
C705 ALU_1b_3/AND_7/out ALU_1b_3/AND_6/w_64_45# 0.13fF
C706 ALU_1b_0/AND_2/out ALU_1b_0/AND_1/a_78_51# 0.24fF
C707 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out vdd 0.06fF
C708 ALU_1b_0/AND_3/out ALU_1b_0/AND_4/out 0.98fF
C709 gnd ALU_1b_3/NOT_5/in 0.07fF
C710 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# vdd 0.22fF
C711 ALU_1b_3/NOR_2/A ALU_1b_3/NOT_4/in 0.03fF
C712 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.05fF
C713 ALU_1b_0/NOR_2/w_n27_1# vdd 0.24fF
C714 ALU_1b_1/decoder_0/AND_3/a_78_51# ALU_1b_1/AND_12/w_64_45# 0.09fF
C715 ALU_1b_2/AND_18/A ALU_1b_2/AND_18/a_78_51# 0.03fF
C716 ALU_1b_1/AND_3/out ALU_1b_1/AND_5/B 0.11fF
C717 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/AND_16/A 0.22fF
C718 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/AND_17/A 0.04fF
C719 ALU_1b_2/full_adder_0/NOR_0/B gnd 0.07fF
C720 S1 ALU_1b_3/decoder_0/AND_3/a_78_51# 0.19fF
C721 gnd ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.04fF
C722 ALU_1b_2/AND_2/a_78_51# B1 0.03fF
C723 ALU_1b_1/AND_19/A ALU_1b_1/NOR_0/A 0.10fF
C724 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/AND_5/out 0.70fF
C725 gnd ALU_1b_2/AND_14/B 0.07fF
C726 vdd ALU_1b_1/decoder_0/AND_0/a_78_51# 0.06fF
C727 ALU_1b_1/decoder_0/AND_2/a_78_51# ALU_1b_1/decoder_0/AND_2/B 0.19fF
C728 ALU_1b_1/AND_17/a_78_51# ALU_1b_1/AND_2/B 0.19fF
C729 ALU_1b_0/AND_18/w_64_45# ALU_1b_0/NOR_3/A 0.03fF
C730 ALU_1b_2/full_adder_1/half_adder_1/A ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C731 vdd ALU_1b_3/comparator_0/w_n220_n67# 0.12fF
C732 ALU_1b_0/full_adder_0/NOR_0/A ALU_1b_0/full_adder_0/NOR_0/B 0.38fF
C733 ALU_1b_2/comparator_0/AND_2/w_64_45# ALU_1b_2/comparator_0/NOR_1/A 0.03fF
C734 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/AND_8/out 0.02fF
C735 ALU_1b_1/AND_3/out gnd 0.11fF
C736 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.09fF
C737 ALU_1b_2/AND_10/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C738 ALU_1b_2/NOR_1/A ALU_1b_2/AND_11/B 0.03fF
C739 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C740 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/AND_7/out 0.05fF
C741 ALU_1b_3/AND_6/out ALU_1b_3/AND_8/out 0.10fF
C742 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# ALU_1b_0/full_adder_0/NOR_0/A 0.03fF
C743 ALU_1b_1/AND_6/out vdd 0.20fF
C744 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/NOR_0/B 0.12fF
C745 A3 ALU_1b_1/AND_9/A 0.31fF
C746 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_2/NOT_1/in 0.03fF
C747 ALU_1b_0/NOR_0/B vdd 0.20fF
C748 ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/A 0.72fF
C749 ALU_1b_0/AND_4/out ALU_1b_0/full_adder_1/NOR_0/B 0.09fF
C750 ALU_1b_1/decoder_0/AND_3/a_78_51# gnd 0.07fF
C751 ALU_1b_2/comparator_0/AND_1/w_64_45# ALU_1b_2/comparator_0/NOR_0/B 0.03fF
C752 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_5/w_64_45# 0.06fF
C753 ALU_1b_0/comparator_0/AND_5/w_64_45# ALU_1b_0/comparator_0/AND_5/a_78_51# 0.09fF
C754 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/AND_7/out 0.61fF
C755 ALU_1b_2/AND_7/w_64_45# ALU_1b_2/AND_9/A 0.39fF
C756 B2 ALU_1b_3/AND_2/B 0.28fF
C757 vdd ALU_1b_3/AND_6/a_78_51# 0.06fF
C758 ALU_1b_0/AND_13/a_78_51# ALU_1b_0/AND_15/A 0.05fF
C759 vdd ALU_1b_2/AND_17/a_78_51# 0.06fF
C760 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_3/A 0.03fF
C761 gnd ALU_1b_3/AND_9/out 0.07fF
C762 ALU_1b_1/AND_3/w_64_45# ALU_1b_1/AND_5/B 0.06fF
C763 ALU_1b_1/comparator_0/AND_5/w_64_45# ALU_1b_1/AND_7/out 0.30fF
C764 vdd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.02fF
C765 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_15/A 0.50fF
C766 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# ALU_1b_0/full_adder_1/NOR_0/B 0.36fF
C767 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/AND_8/out 0.22fF
C768 ALU_1b_1/AND_5/w_64_45# ALU_1b_1/C0 0.10fF
C769 ALU_1b_3/AND_3/out ALU_1b_3/AND_3/a_78_51# 0.05fF
C770 ALU_1b_3/NOR_4/B ALU_1b_3/NOR_4/w_n27_1# 0.09fF
C771 vdd ALU_1b_3/AND_8/w_64_45# 0.14fF
C772 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/w_n39_45# 0.03fF
C773 ALU_1b_0/AND_15/w_64_45# ALU_1b_0/AND_15/A 0.06fF
C774 ALU_1b_0/NOR_3/A gnd 0.23fF
C775 ALU_1b_2/full_adder_0/NOR_0/A vdd 0.03fF
C776 ALU_1b_3/full_adder_1/half_adder_0/w_36_45# ALU_1b_3/AND_3/out 0.09fF
C777 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out 0.09fF
C778 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_0/AND_2/out 0.06fF
C779 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out 0.20fF
C780 ALU_1b_3/AND_1/w_64_45# ALU_1b_3/C0 0.06fF
C781 gnd ALU_1b_3/AND_8/a_78_51# 0.07fF
C782 ALU_1b_0/NOR_1/B ALU_1b_0/NOR_2/A 0.00fF
C783 ALU_1b_1/full_adder_1/w_448_45# ALU_1b_1/full_adder_1/NOR_0/out 0.11fF
C784 ALU_1b_1/AND_19/A ALU_1b_1/NOT_1/w_n36_43# 0.03fF
C785 ALU_1b_0/NOT_5/in ALU_1b_0/NOR_3/A 0.03fF
C786 ALU_1b_1/comparator_0/NOR_2/A vdd 0.03fF
C787 vdd ALU_1b_3/comparator_0/AND_5/a_78_51# 0.06fF
C788 ALU_1b_2/AND_4/out gnd 0.07fF
C789 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_2/full_adder_0/half_adder_1/A 0.03fF
C790 ALU_1b_2/NOR_0/B ALU_1b_2/NOT_2/in 0.15fF
C791 ALU_1b_0/AND_14/B ALU_1b_0/AND_14/a_78_51# 0.19fF
C792 ALU_1b_1/AND_17/A gnd 0.34fF
C793 A0 ALU_1b_0/AND_6/w_64_45# 0.06fF
C794 gnd ALU_1b_3/NOR_1/A 0.51fF
C795 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.52fF
C796 ALU_1b_1/comparator_0/NOR_0/B vdd 0.09fF
C797 ALU_1b_1/comparator_0/w_88_n67# ALU_1b_1/comparator_0/NOR_0/out 0.11fF
C798 F1 ALU_1b_3/AND_9/A 0.28fF
C799 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_74# vdd 0.02fF
C800 ALU_1b_2/AND_3/out ALU_1b_2/AND_4/out 0.98fF
C801 ALU_1b_1/NOR_4/A ALU_1b_1/NOR_1/A 0.01fF
C802 ALU_1b_3/AND_2/w_64_45# ALU_1b_3/AND_2/a_78_51# 0.09fF
C803 ALU_1b_3/AND_3/out ALU_1b_3/AND_4/w_64_45# 0.20fF
C804 ALU_1b_0/comparator_0/w_n195_n67# vdd 0.12fF
C805 ALU_1b_1/comparator_0/NOR_0/out gnd 0.07fF
C806 ALU_1b_3/AND_7/a_78_51# B2 0.19fF
C807 ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/NOR_1/B 0.01fF
C808 ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/comparator_0/NOR_1/a_n14_7# 0.00fF
C809 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C810 ALU_1b_1/AND_2/w_64_45# B3 0.10fF
C811 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/w_36_45# 0.03fF
C812 ALU_1b_3/AND_3/w_64_45# ALU_1b_3/AND_3/a_78_51# 0.09fF
C813 ALU_1b_0/comparator_0/w_n195_n67# ALU_1b_0/comparator_0/NOR_3/A 0.06fF
C814 ALU_1b_0/NOR_0/A ALU_1b_0/AND_5/B 0.01fF
C815 vdd ALU_1b_2/AND_11/a_78_51# 0.06fF
C816 S1 ALU_1b_3/AND_2/B 0.03fF
C817 ALU_1b_0/AND_13/a_78_51# B0 0.19fF
C818 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/AND_11/B 0.10fF
C819 ALU_1b_1/AND_16/a_78_51# vdd 0.06fF
C820 vdd ALU_1b_2/AND_11/B 1.14fF
C821 gnd ALU_1b_2/comparator_0/AND_2/B 0.07fF
C822 ALU_1b_1/AND_18/a_78_51# ALU_1b_1/AND_5/B 0.19fF
C823 A3 ALU_1b_1/AND_3/A 0.03fF
C824 gnd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.02fF
C825 ALU_1b_3/AND_14/w_64_45# B2 0.06fF
C826 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_2/out 0.27fF
C827 ALU_1b_1/full_adder_1/w_448_45# vdd 0.12fF
C828 gnd ALU_1b_2/AND_10/B 0.13fF
C829 vdd ALU_1b_3/comparator_0/w_n39_45# 0.05fF
C830 ALU_1b_1/AND_10/a_78_51# ALU_1b_1/AND_10/B 0.38fF
C831 ALU_1b_2/AND_15/a_78_51# ALU_1b_2/NOR_1/B 0.05fF
C832 ALU_1b_2/full_adder_1/NOR_0/out gnd 0.07fF
C833 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C834 ALU_1b_3/AND_2/out ALU_1b_3/AND_2/w_64_45# 0.03fF
C835 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_6/out 0.05fF
C836 ALU_1b_1/AND_0/a_78_51# gnd 0.07fF
C837 ALU_1b_0/AND_9/A B0 0.28fF
C838 ALU_1b_1/AND_18/w_64_45# vdd 0.15fF
C839 ALU_1b_2/AND_5/w_64_45# ALU_1b_2/AND_5/B 0.06fF
C840 vdd ALU_1b_2/AND_12/w_64_45# 0.47fF
C841 ALU_1b_3/comparator_0/w_n195_n67# ALU_1b_3/comparator_0/NOR_3/out 0.11fF
C842 gnd ALU_1b_2/AND_12/a_78_51# 0.07fF
C843 ALU_1b_1/AND_18/a_78_51# gnd 0.07fF
C844 vdd ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.06fF
C845 ALU_1b_0/comparator_0/NOR_1/A vdd 0.03fF
C846 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_1/AND_16/A 0.13fF
C847 gnd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.11fF
C848 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.00fF
C849 gnd ALU_1b_2/NOR_2/A 0.07fF
C850 ALU_1b_3/decoder_0/AND_1/B ALU_1b_3/AND_2/B 0.17fF
C851 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/NOR_0/A 0.10fF
C852 ALU_1b_1/AND_2/B gnd 0.48fF
C853 ALU_1b_0/AND_16/A ALU_1b_0/AND_16/w_64_45# 0.06fF
C854 ALU_1b_0/comparator_0/w_n220_n67# ALU_1b_0/comparator_0/NOR_2/A 0.06fF
C855 vdd ALU_1b_2/comparator_0/AND_3/a_78_51# 0.06fF
C856 A0 ALU_1b_0/AND_12/a_78_51# 0.19fF
C857 ALU_1b_3/AND_17/w_64_45# ALU_1b_3/AND_17/a_78_51# 0.09fF
C858 ALU_1b_2/AND_4/out F0 0.01fF
C859 F2 ALU_1b_3/NOT_4/in 0.03fF
C860 vdd ALU_1b_2/AND_5/B 0.10fF
C861 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/AND_9/out 0.29fF
C862 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_1/a_78_51# 0.03fF
C863 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.09fF
C864 ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/AND_1/a_78_51# 0.20fF
C865 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_2/a_78_51# 0.19fF
C866 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_5/B 0.17fF
C867 gnd ALU_1b_2/decoder_0/AND_1/a_78_51# 0.07fF
C868 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_9/a_78_51# 0.09fF
C869 ALU_1b_3/AND_9/out ALU_1b_3/AND_10/B 0.06fF
C870 ALU_1b_0/AND_8/out vdd 0.66fF
C871 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_2/full_adder_1/half_adder_1/A 0.03fF
C872 A2 ALU_1b_3/AND_12/w_64_45# 0.18fF
C873 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_5/B 0.05fF
C874 ALU_1b_1/decoder_0/AND_2/B ALU_1b_1/decoder_0/AND_1/B 0.59fF
C875 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C876 vdd ALU_1b_2/comparator_0/w_88_n67# 0.12fF
C877 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/NOR_0/B 0.38fF
C878 ALU_1b_3/AND_3/w_64_45# ALU_1b_3/AND_3/A 0.09fF
C879 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_1/A 0.13fF
C880 S0 ALU_1b_3/AND_12/w_64_45# 0.68fF
C881 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# ALU_1b_2/AND_5/out 0.29fF
C882 ALU_1b_3/NOR_0/B ALU_1b_3/NOR_0/A 0.33fF
C883 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out 0.09fF
C884 ALU_1b_0/NOT_2/in ALU_1b_0/NOR_2/A 0.03fF
C885 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C886 ALU_1b_1/AND_6/out ALU_1b_1/AND_7/out 0.13fF
C887 ALU_1b_1/AND_10/a_78_51# vdd 0.06fF
C888 ALU_1b_0/AND_15/a_78_51# vdd 0.06fF
C889 A2 ALU_1b_3/AND_5/B 0.01fF
C890 ALU_1b_0/NOR_4/B ALU_1b_0/NOR_1/A 0.07fF
C891 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_3/B 0.15fF
C892 ALU_1b_1/comparator_0/NOR_3/A gnd 0.21fF
C893 ALU_1b_0/NOR_0/A ALU_1b_0/NOR_3/A 0.01fF
C894 ALU_1b_2/NOT_3/in ALU_1b_2/NOR_2/w_n27_1# 0.11fF
C895 A1 ALU_1b_2/AND_8/out 0.11fF
C896 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_7/out 0.20fF
C897 ALU_1b_0/AND_9/a_78_51# ALU_1b_0/AND_9/out 0.05fF
C898 ALU_1b_0/AND_7/a_78_51# ALU_1b_0/AND_8/out 0.10fF
C899 vdd ALU_1b_3/AND_3/out 0.03fF
C900 ALU_1b_0/AND_17/A ALU_1b_0/AND_2/B 0.26fF
C901 S0 ALU_1b_3/AND_5/B 0.03fF
C902 ALU_1b_0/comparator_0/w_113_n67# ALU_1b_0/AND_10/B 0.03fF
C903 ALU_1b_1/NOR_4/A ALU_1b_1/NOR_4/w_n27_1# 0.10fF
C904 ALU_1b_2/AND_15/A ALU_1b_2/AND_12/w_64_45# 0.36fF
C905 ALU_1b_2/NOR_0/w_n27_1# ALU_1b_2/NOR_2/A 0.03fF
C906 ALU_1b_3/AND_2/out ALU_1b_3/AND_1/out 0.11fF
C907 C0 ALU_1b_0/AND_5/B 0.01fF
C908 ALU_1b_1/AND_18/a_78_51# ALU_1b_1/NOR_3/A 0.07fF
C909 ALU_1b_3/comparator_0/AND_2/a_78_51# ALU_1b_3/comparator_0/NOR_1/A 0.38fF
C910 ALU_1b_0/AND_4/w_64_45# B0 0.10fF
C911 ALU_1b_1/AND_7/w_64_45# vdd 0.14fF
C912 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C913 ALU_1b_1/comparator_0/NOR_3/out vdd 0.03fF
C914 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_2/AND_5/out 0.04fF
C915 ALU_1b_0/AND_19/w_64_45# vdd 0.15fF
C916 ALU_1b_1/NOT_1/in ALU_1b_1/AND_5/out 0.21fF
C917 ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.10fF
C918 B3 ALU_1b_1/C0 2.32fF
C919 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C920 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out vdd 0.06fF
C921 ALU_1b_0/AND_4/out C1 0.01fF
C922 ALU_1b_1/AND_7/a_78_51# gnd 0.07fF
C923 vdd ALU_1b_3/decoder_0/AND_3/a_78_51# 0.06fF
C924 ALU_1b_0/decoder_0/AND_0/a_78_51# S1 0.02fF
C925 ALU_1b_2/comparator_0/NOR_0/A ALU_1b_2/comparator_0/NOR_0/B 0.33fF
C926 ALU_1b_0/AND_19/a_78_51# gnd 0.07fF
C927 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/w_n39_45# 0.11fF
C928 ALU_1b_2/decoder_0/AND_2/a_78_51# ALU_1b_2/AND_12/w_64_45# 0.09fF
C929 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.10fF
C930 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C931 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_5/a_78_51# 0.29fF
C932 ALU_1b_3/comparator_0/AND_1/a_78_51# ALU_1b_3/comparator_0/NOR_0/B 0.05fF
C933 ALU_1b_2/AND_6/w_64_45# ALU_1b_2/AND_2/B 0.03fF
C934 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/w_448_45# 0.16fF
C935 ALU_1b_1/comparator_0/AND_2/a_78_51# vdd 0.06fF
C936 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_13/a_78_51# 0.09fF
C937 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out 0.14fF
C938 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.09fF
C939 ALU_1b_3/AND_7/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C940 ALU_1b_0/AND_17/A vdd 0.02fF
C941 ALU_1b_3/NOR_1/A ALU_1b_3/NOR_2/A 0.12fF
C942 vdd ALU_1b_3/NOR_0/w_n27_1# 0.12fF
C943 ALU_1b_2/comparator_0/AND_5/a_78_51# ALU_1b_2/AND_7/out 0.14fF
C944 ALU_1b_2/comparator_0/NOR_1/A ALU_1b_2/comparator_0/w_113_n67# 0.06fF
C945 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_74# vdd 0.02fF
C946 ALU_1b_0/AND_8/out ALU_1b_0/comparator_0/AND_4/a_78_51# 0.20fF
C947 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_14/B 0.06fF
C948 ALU_1b_0/AND_15/B ALU_1b_0/AND_15/A 0.28fF
C949 vdd ALU_1b_2/NOR_3/A 0.22fF
C950 ALU_1b_2/decoder_0/AND_2/a_78_51# ALU_1b_2/AND_5/B 0.05fF
C951 gnd ALU_1b_3/AND_15/A 0.87fF
C952 ALU_1b_3/comparator_0/AND_4/w_64_45# ALU_1b_3/AND_8/out 0.37fF
C953 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C954 ALU_1b_0/AND_6/w_64_45# ALU_1b_0/decoder_0/AND_2/B 0.09fF
C955 ALU_1b_1/comparator_0/AND_4/w_64_45# vdd 0.14fF
C956 ALU_1b_3/AND_14/B ALU_1b_3/AND_15/A 0.16fF
C957 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/AND_5/out 0.19fF
C958 ALU_1b_1/AND_15/a_78_51# ALU_1b_1/AND_15/A 0.05fF
C959 ALU_1b_2/NOR_4/w_n27_1# ALU_1b_2/NOR_3/A 0.06fF
C960 vdd ALU_1b_3/AND_3/w_64_45# 0.21fF
C961 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/AND_16/A 0.01fF
C962 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.01fF
C963 ALU_1b_0/full_adder_1/NOR_0/out vdd 0.03fF
C964 ALU_1b_1/AND_18/A ALU_1b_1/AND_5/B 0.26fF
C965 ALU_1b_1/comparator_0/AND_4/a_78_51# gnd 0.07fF
C966 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/A 0.13fF
C967 ALU_1b_0/AND_4/a_78_51# vdd 0.06fF
C968 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_1/A 0.01fF
C969 vdd F1 0.31fF
C970 gnd ALU_1b_3/decoder_0/AND_2/a_78_51# 0.07fF
C971 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C972 ALU_1b_1/full_adder_0/half_adder_1/A gnd 0.03fF
C973 ALU_1b_1/comparator_0/w_113_n67# ALU_1b_1/comparator_0/NOR_1/B 0.62fF
C974 vdd ALU_1b_3/AND_17/A 0.02fF
C975 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C976 ALU_1b_3/NOR_4/A ALU_1b_3/AND_11/a_78_51# 0.07fF
C977 ALU_1b_1/AND_14/a_78_51# ALU_1b_1/AND_15/B 0.05fF
C978 gnd ALU_1b_2/NOT_4/in 0.07fF
C979 ALU_1b_1/AND_19/A ALU_1b_1/AND_5/B 0.26fF
C980 ALU_1b_3/AND_8/w_64_45# ALU_1b_3/C0 0.06fF
C981 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.01fF
C982 ALU_1b_2/AND_1/w_64_45# vdd 0.15fF
C983 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/full_adder_1/half_adder_0/w_36_45# 0.09fF
C984 ALU_1b_0/AND_3/out gnd 0.11fF
C985 ALU_1b_1/AND_18/A gnd 0.27fF
C986 vdd ALU_1b_3/comparator_0/NOR_0/out 0.03fF
C987 ALU_1b_2/AND_7/out ALU_1b_2/comparator_0/w_n39_45# 0.06fF
C988 ALU_1b_1/AND_16/A ALU_1b_1/AND_16/w_64_45# 0.06fF
C989 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_9/out 0.19fF
C990 ALU_1b_0/AND_6/a_78_51# gnd 0.07fF
C991 ALU_1b_3/comparator_0/NOR_0/out ALU_1b_3/comparator_0/NOR_1/B 0.05fF
C992 ALU_1b_0/AND_11/a_78_51# ALU_1b_0/AND_11/B 0.19fF
C993 ALU_1b_2/NOT_6/in ALU_1b_2/NOR_1/A 0.37fF
C994 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/w_36_45# 0.03fF
C995 ALU_1b_0/NOT_1/in ALU_1b_0/AND_18/A 0.12fF
C996 B1 ALU_1b_2/AND_5/B 0.28fF
C997 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_74# vdd 0.02fF
C998 ALU_1b_1/AND_2/a_78_51# vdd 0.06fF
C999 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/w_n195_n67# 0.19fF
C1000 ALU_1b_1/NOR_4/B gnd 0.07fF
C1001 ALU_1b_1/AND_19/A gnd 0.07fF
C1002 ALU_1b_1/AND_8/out B3 0.01fF
C1003 ALU_1b_3/AND_0/out F1 0.01fF
C1004 ALU_1b_0/comparator_0/AND_1/a_78_51# vdd 0.06fF
C1005 ALU_1b_1/comparator_0/NOR_2/out ALU_1b_1/AND_11/B 0.05fF
C1006 ALU_1b_2/AND_16/w_64_45# ALU_1b_2/AND_16/a_78_51# 0.09fF
C1007 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/AND_5/out 0.72fF
C1008 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.03fF
C1009 ALU_1b_0/AND_2/out Cin 0.15fF
C1010 ALU_1b_0/comparator_0/AND_0/w_64_45# ALU_1b_0/comparator_0/NOR_0/A 0.03fF
C1011 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_0/a_78_51# 0.29fF
C1012 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/full_adder_1/half_adder_1/A 0.14fF
C1013 ALU_1b_1/AND_0/w_64_45# ALU_1b_1/AND_0/out 0.09fF
C1014 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# vdd 0.22fF
C1015 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd 0.06fF
C1016 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/AND_4/out 0.20fF
C1017 vdd ALU_1b_3/AND_0/a_78_51# 0.06fF
C1018 ALU_1b_3/AND_17/A ALU_1b_3/full_adder_0/NOR_0/out 0.04fF
C1019 ALU_1b_0/NOT_1/in ALU_1b_0/AND_19/A 0.03fF
C1020 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/AND_5/out 0.05fF
C1021 ALU_1b_1/NOR_0/A vdd 0.20fF
C1022 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_0/half_adder_1/A 0.03fF
C1023 ALU_1b_3/comparator_0/AND_0/w_64_45# ALU_1b_3/comparator_0/AND_2/B 0.06fF
C1024 gnd B2 0.38fF
C1025 ALU_1b_1/AND_6/out ALU_1b_1/AND_9/out 0.29fF
C1026 ALU_1b_0/AND_4/out vdd 0.35fF
C1027 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C1028 ALU_1b_0/NOR_4/A ALU_1b_0/NOT_6/in 0.03fF
C1029 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C1030 ALU_1b_3/AND_14/B B2 0.23fF
C1031 ALU_1b_0/comparator_0/AND_5/w_64_45# vdd 0.13fF
C1032 ALU_1b_1/AND_1/w_64_45# ALU_1b_1/AND_1/out 0.03fF
C1033 vdd ALU_1b_3/AND_18/a_78_51# 0.06fF
C1034 ALU_1b_0/AND_19/w_64_45# ALU_1b_0/AND_19/A 0.06fF
C1035 ALU_1b_3/AND_5/a_78_51# ALU_1b_3/AND_5/B 0.19fF
C1036 ALU_1b_3/decoder_0/AND_2/B ALU_1b_3/AND_12/w_64_45# 0.06fF
C1037 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/w_448_45# 0.06fF
C1038 ALU_1b_0/full_adder_1/NOR_0/B gnd 0.07fF
C1039 ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/AND_2/w_64_45# 0.16fF
C1040 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_5/w_64_45# 0.03fF
C1041 ALU_1b_0/comparator_0/AND_5/a_78_51# gnd 0.07fF
C1042 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.01fF
C1043 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/NOR_1/A 0.03fF
C1044 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/half_adder_1/A 0.14fF
C1045 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/NOR_0/B 0.48fF
C1046 ALU_1b_1/AND_3/out F2 0.01fF
C1047 vdd ALU_1b_3/AND_2/B 0.10fF
C1048 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.09fF
C1049 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# vdd 0.14fF
C1050 ALU_1b_0/NOR_2/A ALU_1b_0/NOT_3/in 0.23fF
C1051 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C1052 ALU_1b_2/AND_0/out ALU_1b_2/AND_2/a_78_51# 0.10fF
C1053 ALU_1b_1/AND_9/A ALU_1b_1/C0 0.28fF
C1054 gnd ALU_1b_2/AND_7/out 0.07fF
C1055 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C1056 ALU_1b_0/AND_14/A vdd 0.03fF
C1057 S1 ALU_1b_1/AND_12/w_64_45# 0.06fF
C1058 ALU_1b_0/AND_19/a_78_51# ALU_1b_0/NOR_0/A 0.16fF
C1059 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/AND_18/A 0.04fF
C1060 ALU_1b_2/AND_2/out ALU_1b_2/AND_1/a_78_51# 0.24fF
C1061 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/NOR_0/A 0.02fF
C1062 ALU_1b_3/AND_0/a_78_51# ALU_1b_3/AND_0/out 0.05fF
C1063 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C1064 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.13fF
C1065 ALU_1b_3/AND_1/a_78_51# ALU_1b_3/AND_2/B 0.19fF
C1066 ALU_1b_3/AND_19/w_64_45# ALU_1b_3/NOR_0/A 0.03fF
C1067 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/full_adder_1/NOR_0/A 0.05fF
C1068 ALU_1b_1/AND_1/w_64_45# ALU_1b_1/C0 0.06fF
C1069 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/AND_16/A 0.01fF
C1070 ALU_1b_0/AND_5/w_64_45# Cin 0.10fF
C1071 ALU_1b_1/AND_7/w_64_45# ALU_1b_1/AND_7/out 0.03fF
C1072 ALU_1b_1/comparator_0/NOR_2/B vdd 0.31fF
C1073 ALU_1b_0/AND_12/w_64_45# ALU_1b_0/AND_5/B 0.03fF
C1074 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.05fF
C1075 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/AND_1/out 0.04fF
C1076 ALU_1b_0/comparator_0/NOR_1/out vdd 0.03fF
C1077 S1 ALU_1b_1/AND_5/B 0.03fF
C1078 ALU_1b_2/AND_2/out ALU_1b_2/AND_0/out 0.96fF
C1079 ALU_1b_1/comparator_0/NOR_2/out gnd 0.07fF
C1080 vdd ALU_1b_3/comparator_0/NOR_3/A 0.03fF
C1081 ALU_1b_2/AND_8/w_64_45# ALU_1b_2/AND_8/a_78_51# 0.09fF
C1082 ALU_1b_3/AND_0/out ALU_1b_3/AND_2/B 0.11fF
C1083 ALU_1b_0/AND_1/w_64_45# ALU_1b_0/AND_1/a_78_51# 0.09fF
C1084 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.03fF
C1085 ALU_1b_2/AND_11/a_78_51# ALU_1b_2/AND_9/A 0.03fF
C1086 ALU_1b_0/AND_3/a_78_51# ALU_1b_0/AND_3/A 0.03fF
C1087 ALU_1b_2/AND_9/A ALU_1b_2/AND_11/B 0.37fF
C1088 ALU_1b_0/full_adder_0/NOR_0/out gnd 0.07fF
C1089 ALU_1b_1/AND_4/out ALU_1b_1/full_adder_1/half_adder_1/A 0.11fF
C1090 ALU_1b_3/AND_9/out ALU_1b_3/AND_7/out 0.02fF
C1091 ALU_1b_3/comparator_0/AND_3/w_64_45# ALU_1b_3/comparator_0/AND_3/a_78_51# 0.09fF
C1092 ALU_1b_0/NOR_2/A ALU_1b_0/NOR_2/w_n27_1# 0.06fF
C1093 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.03fF
C1094 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/AND_1/out 0.06fF
C1095 ALU_1b_1/NOT_1/w_n36_43# vdd 0.06fF
C1096 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out 0.00fF
C1097 ALU_1b_3/AND_12/a_78_51# ALU_1b_3/AND_15/A 0.05fF
C1098 ALU_1b_2/AND_12/w_64_45# ALU_1b_2/decoder_0/AND_1/B 0.03fF
C1099 ALU_1b_0/NOR_3/B vdd 0.33fF
C1100 ALU_1b_1/AND_14/B ALU_1b_1/AND_12/w_64_45# 0.03fF
C1101 S1 gnd 7.53fF
C1102 ALU_1b_2/comparator_0/AND_3/w_64_45# ALU_1b_2/AND_8/out 0.16fF
C1103 ALU_1b_0/decoder_0/AND_2/B S0 0.29fF
C1104 ALU_1b_1/AND_4/a_78_51# B3 0.03fF
C1105 ALU_1b_2/NOT_6/in ALU_1b_2/NOR_4/w_n27_1# 0.11fF
C1106 vdd ALU_1b_3/AND_7/a_78_51# 0.06fF
C1107 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_14/A 0.09fF
C1108 ALU_1b_1/NOR_4/w_n27_1# ALU_1b_1/NOR_3/B 0.20fF
C1109 vdd ALU_1b_2/AND_19/a_78_51# 0.06fF
C1110 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/AND_4/out 0.20fF
C1111 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_0/half_adder_1/A 0.26fF
C1112 ALU_1b_1/comparator_0/AND_4/w_64_45# ALU_1b_1/AND_7/out 0.10fF
C1113 ALU_1b_3/comparator_0/NOR_0/A ALU_1b_3/comparator_0/NOR_0/out 0.03fF
C1114 ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/AND_2/B 0.05fF
C1115 ALU_1b_1/AND_14/A ALU_1b_1/AND_15/A 0.10fF
C1116 ALU_1b_2/full_adder_1/NOR_0/out ALU_1b_2/AND_18/A 0.04fF
C1117 ALU_1b_3/full_adder_0/half_adder_0/w_36_45# ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.09fF
C1118 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.00fF
C1119 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out vdd 0.06fF
C1120 ALU_1b_3/AND_3/out ALU_1b_3/C0 0.01fF
C1121 ALU_1b_2/NOT_5/in gnd 0.07fF
C1122 vdd ALU_1b_3/AND_14/w_64_45# 0.29fF
C1123 ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/w_n39_45# 0.15fF
C1124 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_0/half_adder_1/A 0.03fF
C1125 ALU_1b_1/full_adder_0/NOR_0/B gnd 0.07fF
C1126 S1 ALU_1b_2/decoder_0/AND_3/a_78_51# 0.19fF
C1127 gnd ALU_1b_3/AND_13/a_78_51# 0.07fF
C1128 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out gnd 0.04fF
C1129 ALU_1b_3/AND_13/a_78_51# ALU_1b_3/AND_14/B 0.10fF
C1130 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/w_n74_45# 0.03fF
C1131 ALU_1b_1/AND_8/out ALU_1b_1/AND_9/A 0.12fF
C1132 F1 ALU_1b_3/AND_9/a_78_51# 0.19fF
C1133 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_15/B 0.03fF
C1134 gnd ALU_1b_3/decoder_0/AND_1/B 0.07fF
C1135 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.06fF
C1136 ALU_1b_1/AND_14/B gnd 0.07fF
C1137 vdd ALU_1b_3/comparator_0/AND_4/a_78_51# 0.06fF
C1138 ALU_1b_0/decoder_0/AND_0/a_78_51# vdd 0.06fF
C1139 ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/NOR_0/out 0.15fF
C1140 ALU_1b_0/AND_7/out ALU_1b_0/comparator_0/w_n74_45# 0.10fF
C1141 ALU_1b_2/AND_14/A ALU_1b_2/AND_14/a_78_51# 0.03fF
C1142 ALU_1b_0/AND_15/B ALU_1b_0/AND_15/w_64_45# 0.06fF
C1143 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.09fF
C1144 ALU_1b_1/AND_0/out ALU_1b_1/AND_2/w_64_45# 0.20fF
C1145 ALU_1b_0/NOR_1/B ALU_1b_0/NOR_1/A 0.33fF
C1146 ALU_1b_0/comparator_0/w_n220_n67# ALU_1b_0/comparator_0/NOR_2/B 0.62fF
C1147 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_10/a_78_51# 0.09fF
C1148 ALU_1b_2/AND_3/a_78_51# ALU_1b_2/AND_5/B 0.29fF
C1149 vdd ALU_1b_2/comparator_0/w_n220_n67# 0.12fF
C1150 gnd ALU_1b_3/AND_9/A 0.35fF
C1151 ALU_1b_2/NOT_1/in ALU_1b_2/NOT_1/w_n36_43# 0.06fF
C1152 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.20fF
C1153 ALU_1b_1/AND_15/w_64_45# ALU_1b_1/AND_15/a_78_51# 0.09fF
C1154 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_1/AND_5/out 0.10fF
C1155 ALU_1b_2/AND_16/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.03fF
C1156 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# 0.48fF
C1157 ALU_1b_0/AND_6/out vdd 0.20fF
C1158 ALU_1b_2/comparator_0/w_113_n67# ALU_1b_2/comparator_0/NOR_1/out 0.11fF
C1159 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/A 0.16fF
C1160 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/w_448_45# 0.06fF
C1161 ALU_1b_0/NOR_4/A gnd 0.23fF
C1162 vdd ALU_1b_3/AND_18/A 0.02fF
C1163 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out gnd 0.04fF
C1164 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# ALU_1b_2/full_adder_0/half_adder_1/A 0.06fF
C1165 ALU_1b_3/AND_17/A ALU_1b_3/full_adder_0/w_448_45# 0.03fF
C1166 S1 ALU_1b_3/AND_6/w_64_45# 0.62fF
C1167 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/w_36_45# 0.12fF
C1168 ALU_1b_0/decoder_0/AND_3/a_78_51# gnd 0.07fF
C1169 S1 F0 0.22fF
C1170 ALU_1b_1/AND_2/B F2 0.01fF
C1171 vdd ALU_1b_2/AND_6/a_78_51# 0.06fF
C1172 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOR_4/B 0.09fF
C1173 gnd ALU_1b_3/AND_3/a_78_51# 0.07fF
C1174 ALU_1b_1/AND_17/a_78_51# vdd 0.06fF
C1175 ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# 0.00fF
C1176 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_74# 0.01fF
C1177 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_1/AND_16/A 0.03fF
C1178 ALU_1b_1/comparator_0/AND_0/w_64_45# ALU_1b_1/AND_6/out 0.26fF
C1179 gnd ALU_1b_2/AND_9/out 0.07fF
C1180 ALU_1b_2/AND_16/A ALU_1b_2/AND_16/a_78_51# 0.03fF
C1181 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_2/a_n14_7# 0.00fF
C1182 vdd ALU_1b_3/NOR_4/B 0.03fF
C1183 F1 ALU_1b_3/C0 11.41fF
C1184 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_74# vdd 0.02fF
C1185 vdd ALU_1b_3/AND_19/A 0.03fF
C1186 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/NOR_0/B 0.48fF
C1187 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.05fF
C1188 ALU_1b_0/AND_0/w_64_45# A0 0.10fF
C1189 ALU_1b_0/AND_8/out ALU_1b_0/AND_6/w_64_45# 0.15fF
C1190 ALU_1b_1/AND_4/out ALU_1b_1/AND_5/B 0.38fF
C1191 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/NOR_3/out 0.15fF
C1192 vdd ALU_1b_2/AND_8/w_64_45# 0.14fF
C1193 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_0/out 0.23fF
C1194 ALU_1b_2/AND_4/w_64_45# ALU_1b_2/AND_5/B 0.06fF
C1195 ALU_1b_1/AND_1/out ALU_1b_1/AND_1/a_78_51# 0.05fF
C1196 ALU_1b_1/NOT_3/in ALU_1b_1/NOR_2/B 0.03fF
C1197 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C1198 ALU_1b_0/AND_0/w_64_45# ALU_1b_0/AND_0/a_78_51# 0.09fF
C1199 gnd ALU_1b_2/AND_8/a_78_51# 0.07fF
C1200 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/AND_4/out 0.70fF
C1201 ALU_1b_1/NOT_6/in ALU_1b_1/NOR_4/B 0.15fF
C1202 ALU_1b_1/comparator_0/AND_0/a_78_51# ALU_1b_1/comparator_0/NOR_0/A 0.05fF
C1203 A2 ALU_1b_3/AND_6/a_78_51# 0.19fF
C1204 ALU_1b_0/comparator_0/NOR_2/A vdd 0.03fF
C1205 ALU_1b_0/AND_3/out C0 0.01fF
C1206 ALU_1b_2/AND_17/w_64_45# ALU_1b_2/NOR_3/B 0.07fF
C1207 ALU_1b_3/AND_6/w_64_45# ALU_1b_3/decoder_0/AND_1/B 0.13fF
C1208 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/NOR_0/B 0.05fF
C1209 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.04fF
C1210 Cout vdd 0.12fF
C1211 ALU_1b_0/NOT_4/in ALU_1b_0/NOR_2/w_n27_1# 0.11fF
C1212 C1 gnd 0.31fF
C1213 vdd ALU_1b_2/comparator_0/AND_5/a_78_51# 0.06fF
C1214 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C1215 ALU_1b_1/AND_4/out gnd 0.07fF
C1216 ALU_1b_1/AND_1/out ALU_1b_1/AND_0/out 0.11fF
C1217 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_1/full_adder_1/half_adder_1/A 0.03fF
C1218 ALU_1b_2/AND_3/A ALU_1b_2/AND_5/B 0.42fF
C1219 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.70fF
C1220 ALU_1b_0/AND_0/w_64_45# ALU_1b_0/AND_0/out 0.09fF
C1221 ALU_1b_0/AND_16/a_78_51# ALU_1b_0/AND_2/B 0.19fF
C1222 ALU_1b_1/AND_3/out ALU_1b_1/AND_3/w_64_45# 0.09fF
C1223 ALU_1b_1/AND_19/A ALU_1b_1/AND_19/a_78_51# 0.03fF
C1224 ALU_1b_3/full_adder_1/half_adder_1/w_36_45# ALU_1b_3/full_adder_1/half_adder_1/A 0.06fF
C1225 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C1226 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_5/B 0.16fF
C1227 vdd ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out 0.06fF
C1228 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out 0.05fF
C1229 ALU_1b_3/AND_9/A ALU_1b_3/AND_6/w_64_45# 0.36fF
C1230 Cin B0 2.33fF
C1231 ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/AND_2/a_78_51# 0.03fF
C1232 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_5/a_78_51# 0.05fF
C1233 gnd ALU_1b_2/NOR_1/A 0.51fF
C1234 ALU_1b_3/AND_9/w_64_45# F1 0.06fF
C1235 ALU_1b_3/AND_16/w_64_45# ALU_1b_3/AND_2/B 0.10fF
C1236 ALU_1b_0/comparator_0/NOR_0/B vdd 0.09fF
C1237 ALU_1b_1/AND_10/a_78_51# ALU_1b_1/NOR_1/A 0.05fF
C1238 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C1239 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_1/NOR_0/B 0.00fF
C1240 ALU_1b_3/NOT_1/in ALU_1b_3/AND_18/A 0.12fF
C1241 ALU_1b_0/AND_18/w_64_45# ALU_1b_0/AND_18/a_78_51# 0.09fF
C1242 ALU_1b_1/AND_12/a_78_51# ALU_1b_1/AND_12/w_64_45# 0.09fF
C1243 ALU_1b_2/comparator_0/AND_2/w_64_45# ALU_1b_2/comparator_0/AND_2/a_78_51# 0.09fF
C1244 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_4/w_64_45# 0.03fF
C1245 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/AND_7/out 0.11fF
C1246 ALU_1b_1/AND_1/a_78_51# ALU_1b_1/C0 0.03fF
C1247 ALU_1b_0/comparator_0/NOR_0/out gnd 0.07fF
C1248 ALU_1b_0/AND_8/w_64_45# C0 0.06fF
C1249 ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.26fF
C1250 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C1251 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/NOR_0/out 0.03fF
C1252 ALU_1b_3/NOR_0/B ALU_1b_3/NOR_3/A 0.01fF
C1253 gnd ALU_1b_3/AND_3/A 0.07fF
C1254 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C1255 ALU_1b_1/comparator_0/AND_3/w_64_45# ALU_1b_1/comparator_0/AND_5/B 0.06fF
C1256 ALU_1b_1/NOR_2/B ALU_1b_1/NOR_2/w_n27_1# 0.09fF
C1257 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_2/NOT_1/in 0.03fF
C1258 ALU_1b_1/AND_11/a_78_51# vdd 0.06fF
C1259 S1 ALU_1b_2/AND_2/B 0.03fF
C1260 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_1/AND_5/out 0.04fF
C1261 ALU_1b_3/NOT_1/in ALU_1b_3/AND_19/A 0.03fF
C1262 ALU_1b_0/AND_16/a_78_51# vdd 0.06fF
C1263 vdd ALU_1b_1/AND_11/B 1.14fF
C1264 ALU_1b_0/AND_5/out ALU_1b_0/AND_5/a_78_51# 0.05fF
C1265 ALU_1b_3/NOR_4/A ALU_1b_3/NOT_6/in 0.03fF
C1266 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C1267 ALU_1b_2/NOT_1/in ALU_1b_2/full_adder_1/half_adder_1/A 0.23fF
C1268 ALU_1b_2/AND_2/out ALU_1b_2/C0 0.16fF
C1269 ALU_1b_1/AND_0/out ALU_1b_1/C0 0.01fF
C1270 ALU_1b_1/comparator_0/AND_2/B gnd 0.07fF
C1271 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C1272 ALU_1b_2/AND_7/a_78_51# ALU_1b_2/AND_7/out 0.16fF
C1273 ALU_1b_3/C0 ALU_1b_3/AND_2/B 0.28fF
C1274 S1 ALU_1b_3/decoder_0/AND_1/a_78_51# 0.03fF
C1275 vdd ALU_1b_3/comparator_0/NOR_2/out 0.03fF
C1276 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_4/a_78_8# 0.00fF
C1277 ALU_1b_1/AND_10/B gnd 0.13fF
C1278 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_74# 0.01fF
C1279 vdd ALU_1b_2/comparator_0/w_n39_45# 0.05fF
C1280 ALU_1b_3/full_adder_1/half_adder_0/w_36_45# ALU_1b_3/AND_4/out 0.29fF
C1281 ALU_1b_1/full_adder_1/NOR_0/out gnd 0.07fF
C1282 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_0/NOR_0/B 0.00fF
C1283 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.09fF
C1284 ALU_1b_0/AND_18/w_64_45# vdd 0.15fF
C1285 ALU_1b_3/AND_9/A ALU_1b_3/AND_10/B 0.29fF
C1286 vdd ALU_1b_1/AND_12/w_64_45# 0.47fF
C1287 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.09fF
C1288 ALU_1b_1/AND_12/a_78_51# gnd 0.07fF
C1289 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/w_n74_45# 0.18fF
C1290 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.05fF
C1291 ALU_1b_0/AND_18/a_78_51# gnd 0.07fF
C1292 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out vdd 0.06fF
C1293 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C1294 ALU_1b_2/AND_12/a_78_51# ALU_1b_2/AND_14/B 0.05fF
C1295 ALU_1b_1/NOR_2/A gnd 0.07fF
C1296 ALU_1b_0/AND_0/out ALU_1b_0/AND_2/out 0.96fF
C1297 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_4/a_78_51# 0.04fF
C1298 ALU_1b_3/comparator_0/AND_3/a_78_51# ALU_1b_3/AND_8/out 0.03fF
C1299 ALU_1b_0/AND_2/B gnd 0.48fF
C1300 ALU_1b_3/AND_1/w_64_45# ALU_1b_3/AND_1/out 0.03fF
C1301 ALU_1b_1/comparator_0/AND_3/a_78_51# vdd 0.06fF
C1302 ALU_1b_1/comparator_0/NOR_1/A ALU_1b_1/comparator_0/NOR_1/B 0.33fF
C1303 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_1/A 0.01fF
C1304 ALU_1b_1/AND_13/a_78_51# ALU_1b_1/AND_14/A 0.05fF
C1305 vdd ALU_1b_1/AND_5/B 0.10fF
C1306 ALU_1b_1/AND_4/w_64_45# ALU_1b_1/AND_4/a_78_51# 0.09fF
C1307 ALU_1b_3/decoder_0/AND_1/a_78_51# ALU_1b_3/decoder_0/AND_1/B 0.19fF
C1308 ALU_1b_1/decoder_0/AND_1/a_78_51# gnd 0.07fF
C1309 ALU_1b_2/AND_7/out ALU_1b_2/comparator_0/AND_4/a_78_51# 0.03fF
C1310 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_3/AND_3/out 0.03fF
C1311 ALU_1b_3/AND_4/out ALU_1b_3/AND_4/w_64_45# 0.03fF
C1312 ALU_1b_0/AND_14/A ALU_1b_0/AND_14/B 0.42fF
C1313 ALU_1b_0/AND_9/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C1314 vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.02fF
C1315 ALU_1b_2/NOT_6/in ALU_1b_3/C0 0.03fF
C1316 ALU_1b_2/AND_3/out ALU_1b_2/AND_5/w_64_45# 0.20fF
C1317 ALU_1b_1/comparator_0/w_88_n67# vdd 0.12fF
C1318 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_4/w_n27_1# 0.11fF
C1319 vdd ALU_1b_3/full_adder_0/NOR_0/B 0.91fF
C1320 ALU_1b_3/AND_3/out ALU_1b_3/AND_5/out 0.11fF
C1321 ALU_1b_3/decoder_0/AND_1/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C1322 S0 ALU_1b_2/AND_12/w_64_45# 0.68fF
C1323 vdd gnd 7.21fF
C1324 ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/w_113_n67# 0.02fF
C1325 ALU_1b_2/comparator_0/w_88_n67# ALU_1b_2/comparator_0/NOR_1/B 0.19fF
C1326 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/NOR_0/B 0.38fF
C1327 ALU_1b_0/AND_10/a_78_51# vdd 0.06fF
C1328 vdd ALU_1b_3/AND_14/B 0.03fF
C1329 ALU_1b_0/NOR_0/A ALU_1b_0/NOR_0/w_n27_1# 0.06fF
C1330 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# ALU_1b_2/full_adder_0/NOR_0/B 0.36fF
C1331 ALU_1b_0/comparator_0/NOR_3/A gnd 0.21fF
C1332 gnd ALU_1b_3/comparator_0/NOR_1/B 0.07fF
C1333 ALU_1b_0/AND_19/a_78_51# ALU_1b_0/AND_5/B 0.19fF
C1334 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/AND_1/out 0.10fF
C1335 ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/decoder_0/AND_2/B 0.03fF
C1336 gnd ALU_1b_3/AND_15/B 0.27fF
C1337 ALU_1b_0/comparator_0/w_n220_n67# ALU_1b_0/AND_11/B 0.03fF
C1338 ALU_1b_0/AND_2/out ALU_1b_0/full_adder_0/NOR_0/B 0.09fF
C1339 ALU_1b_2/AND_3/out vdd 0.03fF
C1340 F1 ALU_1b_3/NOR_1/B 0.01fF
C1341 S0 ALU_1b_2/AND_5/B 0.03fF
C1342 ALU_1b_1/AND_15/B ALU_1b_1/AND_15/a_78_51# 0.19fF
C1343 ALU_1b_3/AND_19/w_64_45# ALU_1b_3/AND_5/B 0.06fF
C1344 ALU_1b_1/comparator_0/w_n220_n67# ALU_1b_1/comparator_0/NOR_2/out 0.11fF
C1345 ALU_1b_0/AND_7/w_64_45# vdd 0.14fF
C1346 gnd ALU_1b_3/AND_1/a_78_51# 0.07fF
C1347 ALU_1b_0/comparator_0/NOR_3/out vdd 0.03fF
C1348 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C1349 ALU_1b_0/AND_7/a_78_51# gnd 0.07fF
C1350 ALU_1b_3/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_3/AND_1/out 0.00fF
C1351 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/NOR_3/out 0.03fF
C1352 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/AND_0/out 0.10fF
C1353 vdd ALU_1b_2/decoder_0/AND_3/a_78_51# 0.06fF
C1354 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/NOR_0/out 0.15fF
C1355 ALU_1b_1/AND_16/w_64_45# ALU_1b_1/NOR_0/B 0.03fF
C1356 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C1357 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/NOR_3/B 0.43fF
C1358 gnd ALU_1b_3/AND_0/out 0.11fF
C1359 ALU_1b_3/AND_7/out B2 0.28fF
C1360 ALU_1b_0/comparator_0/AND_2/a_78_51# vdd 0.06fF
C1361 gnd ALU_1b_3/full_adder_0/NOR_0/out 0.07fF
C1362 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_1/half_adder_1/A 0.13fF
C1363 gnd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.11fF
C1364 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/full_adder_0/NOR_0/B 0.00fF
C1365 ALU_1b_0/AND_18/A ALU_1b_0/AND_18/w_64_45# 0.06fF
C1366 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/NOT_1/in 0.06fF
C1367 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_0/a_78_51# 0.14fF
C1368 ALU_1b_2/decoder_0/AND_1/a_78_51# ALU_1b_2/AND_6/w_64_45# 0.09fF
C1369 ALU_1b_0/comparator_0/AND_0/a_78_51# ALU_1b_0/AND_9/out 0.02fF
C1370 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_1/a_78_51# 0.10fF
C1371 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C1372 vdd ALU_1b_2/NOR_0/w_n27_1# 0.12fF
C1373 ALU_1b_0/AND_7/w_64_45# ALU_1b_0/AND_7/a_78_51# 0.09fF
C1374 ALU_1b_1/AND_17/A ALU_1b_1/AND_2/B 0.26fF
C1375 ALU_1b_3/AND_5/out F1 0.01fF
C1376 ALU_1b_0/NOR_1/B B0 0.01fF
C1377 ALU_1b_0/AND_1/out C1 0.01fF
C1378 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out 0.09fF
C1379 ALU_1b_1/NOR_3/A vdd 0.22fF
C1380 ALU_1b_3/comparator_0/AND_0/w_64_45# ALU_1b_3/AND_9/out 0.30fF
C1381 ALU_1b_1/comparator_0/AND_1/w_64_45# ALU_1b_1/comparator_0/AND_1/a_78_51# 0.09fF
C1382 gnd ALU_1b_2/AND_15/A 0.87fF
C1383 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C1384 ALU_1b_0/comparator_0/AND_4/w_64_45# vdd 0.14fF
C1385 ALU_1b_0/AND_2/w_64_45# ALU_1b_0/AND_2/B 0.06fF
C1386 vdd ALU_1b_2/AND_3/w_64_45# 0.21fF
C1387 ALU_1b_3/AND_4/a_78_51# ALU_1b_3/AND_5/B 0.29fF
C1388 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_74# 0.01fF
C1389 S0 ALU_1b_3/decoder_0/AND_3/a_78_51# 0.03fF
C1390 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/half_adder_1/A 0.16fF
C1391 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_2/AND_16/A 0.03fF
C1392 vdd ALU_1b_3/AND_6/w_64_45# 0.48fF
C1393 ALU_1b_0/comparator_0/AND_4/a_78_51# gnd 0.07fF
C1394 ALU_1b_0/AND_3/out ALU_1b_0/AND_5/B 0.11fF
C1395 ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/decoder_0/AND_1/B 0.29fF
C1396 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/w_448_45# 0.06fF
C1397 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_9/A 0.95fF
C1398 A0 ALU_1b_0/AND_15/A 0.42fF
C1399 ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/comparator_0/NOR_2/A 0.03fF
C1400 vdd F0 0.37fF
C1401 vdd ALU_1b_3/AND_4/out 0.35fF
C1402 ALU_1b_3/AND_17/a_78_51# ALU_1b_3/NOR_3/B 0.07fF
C1403 ALU_1b_3/AND_16/A ALU_1b_3/AND_2/B 0.26fF
C1404 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out gnd 0.04fF
C1405 ALU_1b_0/AND_2/a_78_51# ALU_1b_0/AND_2/B 0.29fF
C1406 ALU_1b_0/AND_1/w_64_45# Cin 0.06fF
C1407 gnd ALU_1b_2/decoder_0/AND_2/a_78_51# 0.07fF
C1408 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_2/A 0.33fF
C1409 ALU_1b_2/AND_17/A vdd 0.02fF
C1410 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C1411 ALU_1b_1/NOT_4/in gnd 0.07fF
C1412 ALU_1b_1/AND_2/out ALU_1b_1/AND_1/a_78_51# 0.24fF
C1413 ALU_1b_0/NOR_1/A ALU_1b_0/NOT_3/in 0.03fF
C1414 ALU_1b_2/decoder_0/AND_3/a_78_51# ALU_1b_2/AND_15/A 0.05fF
C1415 ALU_1b_3/NOR_4/w_n27_1# ALU_1b_3/NOR_1/A 0.09fF
C1416 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_4/B 0.03fF
C1417 ALU_1b_3/AND_3/w_64_45# A2 0.10fF
C1418 ALU_1b_0/AND_18/A gnd 0.27fF
C1419 ALU_1b_0/AND_2/w_64_45# vdd 0.15fF
C1420 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_4/a_78_8# 0.00fF
C1421 ALU_1b_0/AND_1/a_78_51# Cin 0.03fF
C1422 vdd ALU_1b_2/comparator_0/NOR_0/out 0.03fF
C1423 ALU_1b_1/AND_0/a_78_51# ALU_1b_1/AND_2/B 0.14fF
C1424 ALU_1b_3/NOT_2/in ALU_1b_3/NOR_0/w_n27_1# 0.11fF
C1425 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_4/a_78_51# 0.18fF
C1426 ALU_1b_1/AND_6/out ALU_1b_1/AND_9/A 0.01fF
C1427 vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.02fF
C1428 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_2/AND_5/out 0.05fF
C1429 ALU_1b_1/AND_2/out ALU_1b_1/AND_0/out 0.96fF
C1430 ALU_1b_0/AND_2/a_78_51# vdd 0.06fF
C1431 vdd ALU_1b_3/comparator_0/AND_2/B 0.03fF
C1432 ALU_1b_2/comparator_0/AND_3/w_64_45# ALU_1b_2/comparator_0/NOR_2/A 0.03fF
C1433 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_3/a_78_51# 0.19fF
C1434 ALU_1b_2/comparator_0/NOR_0/A ALU_1b_2/comparator_0/w_88_n67# 0.06fF
C1435 ALU_1b_0/AND_19/A gnd 0.07fF
C1436 ALU_1b_1/AND_0/w_64_45# A3 0.10fF
C1437 ALU_1b_2/AND_1/w_64_45# ALU_1b_2/AND_1/a_78_51# 0.09fF
C1438 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C1439 C0 C1 6.42fF
C1440 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# ALU_1b_2/full_adder_1/NOR_0/B 0.36fF
C1441 vdd ALU_1b_3/AND_10/B 1.59fF
C1442 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/A 0.06fF
C1443 gnd ALU_1b_3/NOR_2/B 0.07fF
C1444 ALU_1b_0/full_adder_0/half_adder_1/A gnd 0.03fF
C1445 ALU_1b_0/comparator_0/NOR_1/out ALU_1b_0/AND_10/B 0.05fF
C1446 gnd ALU_1b_3/comparator_0/NOR_0/A 0.17fF
C1447 ALU_1b_0/AND_5/w_64_45# ALU_1b_0/AND_5/a_78_51# 0.09fF
C1448 vdd ALU_1b_3/full_adder_1/NOR_0/out 0.03fF
C1449 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/AND_8/out 0.38fF
C1450 ALU_1b_1/NOR_1/B ALU_1b_1/NOT_3/in 0.15fF
C1451 ALU_1b_1/AND_5/out ALU_1b_1/AND_5/a_78_51# 0.05fF
C1452 ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C1453 ALU_1b_2/AND_0/a_78_51# vdd 0.06fF
C1454 ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/AND_10/B 0.09fF
C1455 ALU_1b_0/NOR_0/A vdd 0.20fF
C1456 gnd B1 0.38fF
C1457 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C1458 F3 gnd 0.07fF
C1459 ALU_1b_2/comparator_0/AND_5/w_64_45# ALU_1b_2/AND_8/out 0.32fF
C1460 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_74# vdd 0.02fF
C1461 ALU_1b_2/AND_1/w_64_45# ALU_1b_2/AND_0/out 0.20fF
C1462 ALU_1b_0/comparator_0/AND_4/w_64_45# ALU_1b_0/comparator_0/AND_4/a_78_51# 0.09fF
C1463 ALU_1b_0/AND_7/out ALU_1b_0/AND_8/out 0.40fF
C1464 ALU_1b_2/AND_8/w_64_45# ALU_1b_2/AND_9/A 0.39fF
C1465 vdd ALU_1b_3/AND_12/a_78_51# 0.06fF
C1466 ALU_1b_0/AND_14/a_78_51# ALU_1b_0/AND_15/A 0.00fF
C1467 vdd ALU_1b_2/AND_18/a_78_51# 0.06fF
C1468 ALU_1b_0/NOR_1/A ALU_1b_0/NOR_2/w_n27_1# 0.10fF
C1469 vdd ALU_1b_3/NOR_2/A 0.03fF
C1470 gnd ALU_1b_3/comparator_0/AND_5/B 0.07fF
C1471 ALU_1b_0/AND_6/w_64_45# ALU_1b_0/decoder_0/AND_0/a_78_51# 0.09fF
C1472 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/NOT_1/in 0.06fF
C1473 A0 B0 0.65fF
C1474 ALU_1b_2/AND_3/out B1 0.01fF
C1475 vdd ALU_1b_2/AND_2/B 0.10fF
C1476 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C1477 ALU_1b_1/AND_7/out gnd 0.07fF
C1478 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_1/AND_5/out 0.00fF
C1479 ALU_1b_1/AND_7/w_64_45# B3 0.06fF
C1480 ALU_1b_3/AND_0/a_78_51# A2 0.19fF
C1481 vdd ALU_1b_3/decoder_0/AND_1/a_78_51# 0.06fF
C1482 ALU_1b_2/comparator_0/NOR_1/A ALU_1b_2/comparator_0/NOR_1/out 0.03fF
C1483 ALU_1b_0/AND_1/out vdd 0.35fF
C1484 ALU_1b_0/AND_12/w_64_45# S1 0.06fF
C1485 ALU_1b_0/AND_6/out ALU_1b_0/AND_6/w_64_45# 0.14fF
C1486 gnd ALU_1b_3/AND_9/a_78_51# 0.07fF
C1487 ALU_1b_3/AND_7/out ALU_1b_3/AND_9/A 0.01fF
C1488 ALU_1b_0/full_adder_0/NOR_0/A gnd 0.07fF
C1489 ALU_1b_1/NOR_1/B ALU_1b_1/NOR_2/w_n27_1# 0.06fF
C1490 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C1491 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_2/full_adder_1/half_adder_1/A 0.26fF
C1492 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_6/w_64_45# 0.09fF
C1493 ALU_1b_3/AND_3/out ALU_1b_3/AND_5/a_78_51# 0.10fF
C1494 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C1495 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_74# 0.01fF
C1496 ALU_1b_0/comparator_0/NOR_2/B vdd 0.31fF
C1497 ALU_1b_0/AND_0/out B0 0.01fF
C1498 A2 ALU_1b_3/AND_2/B 0.50fF
C1499 ALU_1b_2/NOR_0/A ALU_1b_2/NOT_2/in 0.03fF
C1500 ALU_1b_0/AND_15/w_64_45# ALU_1b_0/NOR_1/B 0.06fF
C1501 ALU_1b_0/AND_5/B S1 0.03fF
C1502 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# ALU_1b_1/full_adder_0/half_adder_1/A 0.06fF
C1503 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/w_448_45# 0.16fF
C1504 ALU_1b_0/comparator_0/NOR_2/out gnd 0.07fF
C1505 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_11/a_78_51# 0.09fF
C1506 ALU_1b_3/NOT_1/in ALU_1b_3/full_adder_1/NOR_0/out 0.10fF
C1507 vdd ALU_1b_2/comparator_0/NOR_3/A 0.03fF
C1508 ALU_1b_1/full_adder_0/NOR_0/A vdd 0.03fF
C1509 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_11/B 0.11fF
C1510 ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/comparator_0/NOR_1/out 0.25fF
C1511 C0 ALU_1b_0/AND_2/B 0.01fF
C1512 ALU_1b_2/C0 ALU_1b_2/AND_5/B 0.28fF
C1513 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C1514 vdd ALU_1b_3/full_adder_0/half_adder_1/w_36_45# 0.14fF
C1515 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_16/A 0.23fF
C1516 ALU_1b_1/comparator_0/w_n195_n67# ALU_1b_1/comparator_0/NOR_3/B 0.06fF
C1517 ALU_1b_3/AND_17/A ALU_1b_3/AND_17/w_64_45# 0.06fF
C1518 ALU_1b_0/NOT_1/w_n36_43# vdd 0.06fF
C1519 ALU_1b_2/NOR_4/B ALU_1b_2/NOR_1/A 0.07fF
C1520 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C1521 ALU_1b_1/full_adder_1/NOR_0/A gnd 0.07fF
C1522 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_0/NOT_1/in 0.03fF
C1523 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/AND_5/out 0.70fF
C1524 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/A 0.16fF
C1525 ALU_1b_0/NOR_4/A ALU_1b_0/AND_11/a_78_51# 0.07fF
C1526 ALU_1b_0/comparator_0/AND_0/w_64_45# ALU_1b_0/comparator_0/AND_0/a_78_51# 0.09fF
C1527 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_2/B 0.40fF
C1528 ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.13fF
C1529 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/AND_5/out 0.08fF
C1530 vdd ALU_1b_2/AND_7/a_78_51# 0.06fF
C1531 ALU_1b_1/AND_19/a_78_51# vdd 0.06fF
C1532 ALU_1b_1/AND_4/out F2 0.01fF
C1533 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_1/w_64_45# 0.10fF
C1534 gnd ALU_1b_3/C0 0.53fF
C1535 ALU_1b_1/AND_1/out ALU_1b_1/AND_16/A 0.11fF
C1536 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_3/out 0.05fF
C1537 C0 vdd 0.25fF
C1538 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# ALU_1b_1/AND_0/out 0.09fF
C1539 ALU_1b_2/AND_16/a_78_51# ALU_1b_2/NOR_0/B 0.05fF
C1540 ALU_1b_0/NOT_1/in ALU_1b_0/AND_5/out 0.21fF
C1541 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_1/NOR_0/A 0.06fF
C1542 ALU_1b_2/full_adder_0/half_adder_0/w_36_45# ALU_1b_2/full_adder_0/NOR_0/B 0.12fF
C1543 ALU_1b_2/AND_7/out ALU_1b_2/AND_6/w_64_45# 0.13fF
C1544 ALU_1b_1/NOT_5/in gnd 0.07fF
C1545 vdd ALU_1b_2/AND_14/w_64_45# 0.29fF
C1546 ALU_1b_3/AND_0/w_64_45# ALU_1b_3/AND_0/a_78_51# 0.09fF
C1547 ALU_1b_2/NOR_2/A ALU_1b_2/NOT_4/in 0.03fF
C1548 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.05fF
C1549 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C1550 ALU_1b_0/decoder_0/AND_3/a_78_51# ALU_1b_0/AND_12/w_64_45# 0.09fF
C1551 ALU_1b_1/AND_18/A ALU_1b_1/AND_18/a_78_51# 0.03fF
C1552 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/AND_16/A 0.22fF
C1553 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out 0.05fF
C1554 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/NOR_0/A 0.12fF
C1555 ALU_1b_1/decoder_0/AND_3/a_78_51# S1 0.19fF
C1556 gnd ALU_1b_2/AND_13/a_78_51# 0.07fF
C1557 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out gnd 0.04fF
C1558 ALU_1b_1/AND_2/a_78_51# B3 0.03fF
C1559 ALU_1b_0/AND_19/A ALU_1b_0/NOR_0/A 0.10fF
C1560 gnd ALU_1b_2/decoder_0/AND_1/B 0.07fF
C1561 ALU_1b_0/AND_14/B gnd 0.07fF
C1562 ALU_1b_3/AND_0/w_64_45# ALU_1b_3/AND_2/B 0.06fF
C1563 ALU_1b_0/decoder_0/AND_2/a_78_51# ALU_1b_0/decoder_0/AND_2/B 0.19fF
C1564 vdd ALU_1b_2/comparator_0/AND_4/a_78_51# 0.06fF
C1565 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/NOR_0/B 0.00fF
C1566 ALU_1b_3/AND_19/w_64_45# ALU_1b_3/AND_19/a_78_51# 0.09fF
C1567 ALU_1b_0/AND_17/a_78_51# ALU_1b_0/AND_2/B 0.19fF
C1568 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.01fF
C1569 ALU_1b_1/full_adder_1/half_adder_1/A ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C1570 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# ALU_1b_1/AND_5/out 0.29fF
C1571 ALU_1b_1/comparator_0/w_n220_n67# vdd 0.12fF
C1572 ALU_1b_1/comparator_0/AND_2/w_64_45# ALU_1b_1/comparator_0/NOR_1/A 0.03fF
C1573 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/AND_8/out 0.02fF
C1574 ALU_1b_1/NOR_1/B ALU_1b_1/C0 0.01fF
C1575 gnd ALU_1b_2/AND_9/A 0.35fF
C1576 ALU_1b_1/AND_10/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C1577 ALU_1b_3/AND_17/w_64_45# ALU_1b_3/AND_2/B 0.06fF
C1578 ALU_1b_1/NOR_1/A ALU_1b_1/AND_11/B 0.03fF
C1579 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_2/full_adder_1/half_adder_1/A 0.03fF
C1580 ALU_1b_3/NOR_2/A ALU_1b_3/NOR_2/B 0.47fF
C1581 ALU_1b_1/NOR_4/A ALU_1b_1/AND_9/w_64_45# 0.03fF
C1582 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/AND_16/A 0.06fF
C1583 ALU_1b_2/AND_6/out ALU_1b_2/AND_8/out 0.10fF
C1584 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/AND_7/out 0.05fF
C1585 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C1586 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/NOR_0/B 0.12fF
C1587 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_3/NOT_1/in 0.03fF
C1588 ALU_1b_3/AND_2/out ALU_1b_3/AND_2/a_78_51# 0.05fF
C1589 ALU_1b_0/full_adder_1/NOR_0/A ALU_1b_0/full_adder_1/w_448_45# 0.06fF
C1590 A0 ALU_1b_0/AND_9/A 0.31fF
C1591 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_1/NOT_1/in 0.03fF
C1592 vdd ALU_1b_2/AND_18/A 0.02fF
C1593 ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/A 0.72fF
C1594 ALU_1b_3/NOR_3/B ALU_1b_3/NOR_3/A 0.34fF
C1595 gnd ALU_1b_3/comparator_0/NOR_3/B 0.21fF
C1596 S1 ALU_1b_2/AND_6/w_64_45# 0.62fF
C1597 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_1/out 0.72fF
C1598 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.03fF
C1599 ALU_1b_1/comparator_0/AND_1/w_64_45# ALU_1b_1/comparator_0/NOR_0/B 0.03fF
C1600 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_5/w_64_45# 0.06fF
C1601 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_8/out 0.11fF
C1602 ALU_1b_1/AND_6/a_78_51# vdd 0.06fF
C1603 ALU_1b_1/AND_7/w_64_45# ALU_1b_1/AND_9/A 0.39fF
C1604 B1 ALU_1b_2/AND_2/B 0.28fF
C1605 gnd ALU_1b_2/AND_3/a_78_51# 0.07fF
C1606 ALU_1b_0/AND_17/a_78_51# vdd 0.06fF
C1607 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_3/A 0.03fF
C1608 ALU_1b_1/AND_9/out gnd 0.07fF
C1609 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# vdd 0.14fF
C1610 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.00fF
C1611 vdd ALU_1b_2/NOR_4/B 0.03fF
C1612 ALU_1b_0/comparator_0/AND_5/w_64_45# ALU_1b_0/AND_7/out 0.30fF
C1613 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_15/A 0.50fF
C1614 ALU_1b_3/AND_4/out ALU_1b_3/C0 0.16fF
C1615 ALU_1b_0/AND_8/a_78_51# ALU_1b_0/AND_8/out 0.22fF
C1616 vdd ALU_1b_2/AND_19/A 0.03fF
C1617 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# 0.03fF
C1618 ALU_1b_2/AND_3/out ALU_1b_2/AND_3/a_78_51# 0.05fF
C1619 C1 ALU_1b_0/AND_5/B 0.01fF
C1620 ALU_1b_1/AND_5/out ALU_1b_1/C0 0.01fF
C1621 ALU_1b_2/NOR_4/B ALU_1b_2/NOR_4/w_n27_1# 0.09fF
C1622 ALU_1b_3/AND_8/w_64_45# ALU_1b_3/AND_8/out 0.03fF
C1623 ALU_1b_3/AND_9/out ALU_1b_3/AND_9/A 0.04fF
C1624 ALU_1b_3/comparator_0/AND_3/a_78_51# ALU_1b_3/comparator_0/NOR_2/A 0.17fF
C1625 ALU_1b_1/AND_8/w_64_45# vdd 0.14fF
C1626 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/w_n39_45# 0.03fF
C1627 gnd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.14fF
C1628 ALU_1b_2/full_adder_1/half_adder_0/w_36_45# ALU_1b_2/AND_3/out 0.09fF
C1629 ALU_1b_2/AND_1/w_64_45# ALU_1b_2/C0 0.06fF
C1630 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/AND_5/out 0.20fF
C1631 ALU_1b_1/AND_8/a_78_51# gnd 0.07fF
C1632 vdd F2 0.37fF
C1633 ALU_1b_0/AND_19/A ALU_1b_0/NOT_1/w_n36_43# 0.03fF
C1634 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_1/NOR_0/B 0.00fF
C1635 ALU_1b_3/comparator_0/AND_5/a_78_51# ALU_1b_3/AND_8/out 0.02fF
C1636 ALU_1b_1/comparator_0/AND_5/a_78_51# vdd 0.06fF
C1637 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_14/a_78_51# 0.09fF
C1638 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C1639 ALU_1b_1/NOR_0/B ALU_1b_1/NOT_2/in 0.15fF
C1640 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/NOR_0/A 0.04fF
C1641 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# ALU_1b_0/AND_3/out 0.09fF
C1642 Cout ALU_1b_1/NOR_4/w_n27_1# 0.03fF
C1643 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out vdd 0.06fF
C1644 ALU_1b_3/full_adder_1/NOR_0/A gnd 0.07fF
C1645 ALU_1b_1/NOR_1/A gnd 0.51fF
C1646 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.52fF
C1647 vdd ALU_1b_3/AND_7/out 0.34fF
C1648 ALU_1b_0/comparator_0/w_88_n67# ALU_1b_0/comparator_0/NOR_0/out 0.11fF
C1649 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C1650 F0 ALU_1b_2/AND_9/A 0.28fF
C1651 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# ALU_1b_1/full_adder_0/NOR_0/B 0.36fF
C1652 ALU_1b_1/AND_3/out ALU_1b_1/AND_4/out 0.98fF
C1653 ALU_1b_2/AND_2/w_64_45# ALU_1b_2/AND_2/a_78_51# 0.09fF
C1654 ALU_1b_3/comparator_0/w_88_n67# ALU_1b_3/comparator_0/NOR_0/B 0.20fF
C1655 ALU_1b_2/AND_3/out ALU_1b_2/AND_4/w_64_45# 0.20fF
C1656 ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/NOR_1/B 0.01fF
C1657 ALU_1b_2/AND_7/a_78_51# B1 0.19fF
C1658 ALU_1b_3/NOR_0/B ALU_1b_3/NOR_0/w_n27_1# 0.06fF
C1659 ALU_1b_0/AND_5/out ALU_1b_0/AND_4/out 0.11fF
C1660 ALU_1b_3/NOR_1/A ALU_1b_3/AND_9/A 0.03fF
C1661 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_3/AND_16/A 0.03fF
C1662 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/AND_16/A 0.05fF
C1663 ALU_1b_2/AND_3/w_64_45# ALU_1b_2/AND_3/a_78_51# 0.09fF
C1664 gnd ALU_1b_2/AND_3/A 0.07fF
C1665 ALU_1b_0/AND_1/w_64_45# ALU_1b_0/AND_0/out 0.20fF
C1666 ALU_1b_0/AND_11/a_78_51# vdd 0.06fF
C1667 S1 ALU_1b_1/AND_2/B 0.03fF
C1668 ALU_1b_0/AND_11/B vdd 1.14fF
C1669 gnd ALU_1b_3/AND_16/A 0.14fF
C1670 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# ALU_1b_0/AND_5/out 0.29fF
C1671 ALU_1b_0/comparator_0/AND_2/B gnd 0.07fF
C1672 ALU_1b_0/AND_18/a_78_51# ALU_1b_0/AND_5/B 0.19fF
C1673 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C1674 A0 ALU_1b_0/AND_3/A 0.03fF
C1675 ALU_1b_2/AND_14/w_64_45# B1 0.06fF
C1676 gnd ALU_1b_3/NOR_1/B 0.22fF
C1677 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/NOR_2/out 0.27fF
C1678 ALU_1b_0/AND_10/B gnd 0.13fF
C1679 vdd ALU_1b_2/comparator_0/NOR_2/out 0.03fF
C1680 S1 ALU_1b_2/decoder_0/AND_1/a_78_51# 0.03fF
C1681 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out 0.09fF
C1682 ALU_1b_0/AND_0/out ALU_1b_0/AND_1/a_78_51# 0.10fF
C1683 vdd ALU_1b_1/comparator_0/w_n39_45# 0.05fF
C1684 ALU_1b_0/AND_10/a_78_51# ALU_1b_0/AND_10/B 0.38fF
C1685 ALU_1b_1/AND_15/a_78_51# ALU_1b_1/NOR_1/B 0.05fF
C1686 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# 0.09fF
C1687 ALU_1b_3/AND_18/w_64_45# ALU_1b_3/AND_5/B 0.10fF
C1688 ALU_1b_2/AND_2/out ALU_1b_2/AND_2/w_64_45# 0.03fF
C1689 gnd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_36# 0.02fF
C1690 ALU_1b_3/AND_15/A B2 0.28fF
C1691 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# ALU_1b_0/full_adder_1/NOR_0/B 0.12fF
C1692 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_10/B 0.20fF
C1693 ALU_1b_3/AND_1/out F1 0.01fF
C1694 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/AND_2/out 0.20fF
C1695 ALU_1b_1/AND_5/w_64_45# ALU_1b_1/AND_5/B 0.06fF
C1696 ALU_1b_3/AND_2/w_64_45# ALU_1b_3/AND_2/B 0.06fF
C1697 ALU_1b_0/AND_12/w_64_45# vdd 0.47fF
C1698 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_1/A 0.13fF
C1699 ALU_1b_2/comparator_0/w_n195_n67# ALU_1b_2/comparator_0/NOR_3/out 0.11fF
C1700 ALU_1b_0/AND_12/a_78_51# gnd 0.07fF
C1701 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.09fF
C1702 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C1703 ALU_1b_0/NOR_2/A gnd 0.07fF
C1704 ALU_1b_3/NOT_4/in ALU_1b_3/NOR_2/B 0.15fF
C1705 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/AND_5/out 0.19fF
C1706 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/NOR_0/A 0.10fF
C1707 gnd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# 0.02fF
C1708 ALU_1b_2/decoder_0/AND_1/B ALU_1b_2/AND_2/B 0.17fF
C1709 ALU_1b_0/comparator_0/AND_3/a_78_51# vdd 0.06fF
C1710 ALU_1b_2/AND_17/w_64_45# ALU_1b_2/AND_17/a_78_51# 0.09fF
C1711 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.09fF
C1712 ALU_1b_0/AND_5/B vdd 0.10fF
C1713 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_1/a_78_51# 0.03fF
C1714 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/AND_9/out 0.29fF
C1715 ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/AND_1/a_78_51# 0.20fF
C1716 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/AND_2/a_78_51# 0.19fF
C1717 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_5/B 0.17fF
C1718 ALU_1b_0/decoder_0/AND_1/a_78_51# gnd 0.07fF
C1719 gnd ALU_1b_3/AND_5/out 0.62fF
C1720 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_9/a_78_51# 0.09fF
C1721 ALU_1b_2/AND_9/out ALU_1b_2/AND_10/B 0.06fF
C1722 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_1/full_adder_1/half_adder_1/A 0.03fF
C1723 A1 ALU_1b_2/AND_12/w_64_45# 0.18fF
C1724 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_2/w_64_45# 0.06fF
C1725 ALU_1b_3/comparator_0/AND_1/w_64_45# ALU_1b_3/AND_9/out 0.39fF
C1726 vdd ALU_1b_3/full_adder_0/half_adder_0/w_36_45# 0.14fF
C1727 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_5/B 0.05fF
C1728 vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.02fF
C1729 ALU_1b_0/decoder_0/AND_2/B ALU_1b_0/decoder_0/AND_1/B 0.59fF
C1730 ALU_1b_0/comparator_0/w_88_n67# vdd 0.12fF
C1731 ALU_1b_2/full_adder_0/NOR_0/B vdd 0.91fF
C1732 ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/NOR_0/B 0.10fF
C1733 ALU_1b_2/AND_3/w_64_45# ALU_1b_2/AND_3/A 0.09fF
C1734 ALU_1b_1/AND_12/w_64_45# S0 0.68fF
C1735 vdd ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.06fF
C1736 ALU_1b_2/NOR_0/B ALU_1b_2/NOR_0/A 0.33fF
C1737 ALU_1b_0/AND_6/out ALU_1b_0/AND_7/out 0.13fF
C1738 vdd ALU_1b_2/AND_14/B 0.03fF
C1739 A1 ALU_1b_2/AND_5/B 0.01fF
C1740 gnd ALU_1b_2/comparator_0/NOR_1/B 0.07fF
C1741 ALU_1b_1/NOT_3/in ALU_1b_1/NOR_2/w_n27_1# 0.11fF
C1742 A3 ALU_1b_1/AND_8/out 0.11fF
C1743 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_7/out 0.20fF
C1744 gnd ALU_1b_2/AND_15/B 0.27fF
C1745 ALU_1b_1/AND_3/out vdd 0.03fF
C1746 S0 ALU_1b_1/AND_5/B 0.03fF
C1747 ALU_1b_1/AND_15/A ALU_1b_1/AND_12/w_64_45# 0.36fF
C1748 ALU_1b_1/NOR_0/w_n27_1# ALU_1b_1/NOR_2/A 0.03fF
C1749 ALU_1b_2/AND_2/out ALU_1b_2/AND_1/out 0.11fF
C1750 ALU_1b_0/AND_18/a_78_51# ALU_1b_0/NOR_3/A 0.07fF
C1751 ALU_1b_2/AND_1/a_78_51# gnd 0.07fF
C1752 ALU_1b_2/comparator_0/AND_2/a_78_51# ALU_1b_2/comparator_0/NOR_1/A 0.38fF
C1753 ALU_1b_3/NOR_4/A ALU_1b_3/NOR_4/B 0.35fF
C1754 ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C1755 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.01fF
C1756 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_1/AND_5/out 0.04fF
C1757 ALU_1b_3/AND_18/w_64_45# ALU_1b_3/NOR_3/A 0.03fF
C1758 ALU_1b_3/full_adder_0/half_adder_0/w_36_45# ALU_1b_3/AND_0/out 0.09fF
C1759 gnd A2 0.48fF
C1760 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/NOR_0/out 0.03fF
C1761 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/full_adder_0/w_448_45# 0.11fF
C1762 ALU_1b_1/comparator_0/NOR_0/A ALU_1b_1/comparator_0/NOR_0/B 0.33fF
C1763 ALU_1b_1/decoder_0/AND_3/a_78_51# vdd 0.06fF
C1764 ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.14fF
C1765 ALU_1b_1/decoder_0/AND_2/a_78_51# ALU_1b_1/AND_12/w_64_45# 0.09fF
C1766 S0 gnd 0.48fF
C1767 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.10fF
C1768 ALU_1b_2/AND_0/out gnd 0.11fF
C1769 ALU_1b_1/AND_6/w_64_45# ALU_1b_1/AND_2/B 0.03fF
C1770 S1 ALU_1b_3/decoder_0/AND_2/a_78_51# 0.02fF
C1771 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/w_448_45# 0.16fF
C1772 ALU_1b_2/comparator_0/AND_1/a_78_51# ALU_1b_2/comparator_0/NOR_0/B 0.05fF
C1773 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_5/a_78_51# 0.29fF
C1774 vdd ALU_1b_3/AND_9/out 0.86fF
C1775 ALU_1b_2/full_adder_0/NOR_0/out gnd 0.07fF
C1776 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_13/a_78_51# 0.09fF
C1777 ALU_1b_2/AND_7/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C1778 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C1779 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/AND_2/out 0.70fF
C1780 ALU_1b_2/NOR_1/A ALU_1b_2/NOR_2/A 0.12fF
C1781 gnd ALU_1b_3/NOT_2/in 0.07fF
C1782 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/AND_7/out 0.61fF
C1783 ALU_1b_3/comparator_0/AND_5/w_64_45# ALU_1b_3/comparator_0/AND_5/a_78_51# 0.09fF
C1784 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C1785 ALU_1b_1/comparator_0/AND_5/a_78_51# ALU_1b_1/AND_7/out 0.14fF
C1786 ALU_1b_1/comparator_0/NOR_1/A ALU_1b_1/comparator_0/w_113_n67# 0.06fF
C1787 ALU_1b_1/NOR_0/w_n27_1# vdd 0.12fF
C1788 ALU_1b_3/AND_13/a_78_51# ALU_1b_3/AND_15/A 0.05fF
C1789 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_14/B 0.06fF
C1790 ALU_1b_3/AND_4/out ALU_1b_3/AND_5/out 0.11fF
C1791 ALU_1b_0/NOR_3/A vdd 0.22fF
C1792 ALU_1b_1/AND_5/a_78_51# ALU_1b_1/C0 0.03fF
C1793 ALU_1b_1/decoder_0/AND_2/a_78_51# ALU_1b_1/AND_5/B 0.05fF
C1794 ALU_1b_1/AND_15/A gnd 0.87fF
C1795 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/AND_5/out 0.70fF
C1796 ALU_1b_2/comparator_0/AND_4/w_64_45# ALU_1b_2/AND_8/out 0.37fF
C1797 ALU_1b_2/AND_14/B ALU_1b_2/AND_15/A 0.16fF
C1798 vdd ALU_1b_3/AND_8/a_78_51# 0.06fF
C1799 ALU_1b_0/AND_15/a_78_51# ALU_1b_0/AND_15/A 0.05fF
C1800 ALU_1b_1/NOR_4/w_n27_1# ALU_1b_1/NOR_3/A 0.06fF
C1801 ALU_1b_1/AND_3/w_64_45# vdd 0.21fF
C1802 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/AND_16/A 0.01fF
C1803 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_0/full_adder_0/NOR_0/B 0.00fF
C1804 vdd ALU_1b_2/AND_6/w_64_45# 0.48fF
C1805 S0 ALU_1b_2/decoder_0/AND_3/a_78_51# 0.03fF
C1806 ALU_1b_0/AND_18/A ALU_1b_0/AND_5/B 0.26fF
C1807 ALU_1b_3/AND_15/w_64_45# ALU_1b_3/AND_15/A 0.06fF
C1808 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_1/A 0.01fF
C1809 vdd ALU_1b_2/AND_4/out 0.35fF
C1810 ALU_1b_0/NOT_6/in ALU_1b_2/C0 0.03fF
C1811 ALU_1b_3/NOR_1/B ALU_1b_3/NOR_2/A 0.00fF
C1812 ALU_1b_1/decoder_0/AND_2/a_78_51# gnd 0.07fF
C1813 ALU_1b_0/comparator_0/w_113_n67# ALU_1b_0/comparator_0/NOR_1/B 0.62fF
C1814 ALU_1b_1/AND_17/A vdd 0.02fF
C1815 vdd ALU_1b_3/NOR_1/A 0.22fF
C1816 ALU_1b_2/NOR_4/A ALU_1b_2/AND_11/a_78_51# 0.07fF
C1817 ALU_1b_0/AND_14/a_78_51# ALU_1b_0/AND_15/B 0.05fF
C1818 ALU_1b_0/NOT_4/in gnd 0.07fF
C1819 ALU_1b_0/AND_19/A ALU_1b_0/AND_5/B 0.26fF
C1820 ALU_1b_2/AND_8/w_64_45# ALU_1b_2/C0 0.06fF
C1821 gnd ALU_1b_3/AND_14/a_78_51# 0.07fF
C1822 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/full_adder_1/half_adder_0/w_36_45# 0.09fF
C1823 vdd ALU_1b_1/comparator_0/NOR_0/out 0.03fF
C1824 ALU_1b_1/AND_7/out ALU_1b_1/comparator_0/w_n39_45# 0.06fF
C1825 ALU_1b_3/AND_14/B ALU_1b_3/AND_14/a_78_51# 0.19fF
C1826 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# vdd 0.14fF
C1827 A2 ALU_1b_3/AND_6/w_64_45# 0.06fF
C1828 ALU_1b_3/AND_3/out ALU_1b_3/AND_4/a_78_51# 0.10fF
C1829 vdd ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.02fF
C1830 ALU_1b_2/comparator_0/NOR_0/out ALU_1b_2/comparator_0/NOR_1/B 0.05fF
C1831 ALU_1b_1/NOT_6/in ALU_1b_1/NOR_1/A 0.37fF
C1832 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.01fF
C1833 B3 ALU_1b_1/AND_5/B 0.28fF
C1834 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/NOR_0/B 0.48fF
C1835 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/w_n195_n67# 0.19fF
C1836 S0 F0 0.22fF
C1837 vdd ALU_1b_2/comparator_0/AND_2/B 0.03fF
C1838 ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/comparator_0/NOR_1/a_n14_7# 0.00fF
C1839 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/AND_3/out 0.10fF
C1840 ALU_1b_0/AND_8/out B0 0.01fF
C1841 ALU_1b_2/AND_0/out F0 0.01fF
C1842 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_3/AND_1/out 0.04fF
C1843 ALU_1b_0/comparator_0/NOR_2/out ALU_1b_0/AND_11/B 0.05fF
C1844 ALU_1b_1/AND_16/w_64_45# ALU_1b_1/AND_16/a_78_51# 0.09fF
C1845 vdd ALU_1b_2/AND_10/B 1.59fF
C1846 ALU_1b_3/comparator_0/w_n195_n67# ALU_1b_3/comparator_0/NOR_3/A 0.06fF
C1847 gnd ALU_1b_2/NOR_2/B 0.07fF
C1848 ALU_1b_3/NOR_0/A ALU_1b_3/AND_5/B 0.01fF
C1849 gnd ALU_1b_2/comparator_0/NOR_0/A 0.17fF
C1850 vdd ALU_1b_2/full_adder_1/NOR_0/out 0.03fF
C1851 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/AND_11/B 0.10fF
C1852 ALU_1b_3/AND_13/a_78_51# B2 0.19fF
C1853 ALU_1b_2/AND_17/A ALU_1b_2/full_adder_0/NOR_0/out 0.04fF
C1854 ALU_1b_1/AND_0/a_78_51# vdd 0.06fF
C1855 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/AND_5/out 0.05fF
C1856 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_0/half_adder_1/A 0.03fF
C1857 ALU_1b_2/comparator_0/AND_0/w_64_45# ALU_1b_2/comparator_0/AND_2/B 0.06fF
C1858 ALU_1b_0/AND_6/out ALU_1b_0/AND_9/out 0.29fF
C1859 B3 gnd 0.38fF
C1860 vdd ALU_1b_2/AND_12/a_78_51# 0.06fF
C1861 ALU_1b_2/AND_14/B B1 0.23fF
C1862 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/AND_1/out 0.72fF
C1863 ALU_1b_0/NOR_1/B Cin 0.01fF
C1864 ALU_1b_1/AND_18/a_78_51# vdd 0.06fF
C1865 vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C1866 ALU_1b_2/AND_5/a_78_51# ALU_1b_2/AND_5/B 0.19fF
C1867 ALU_1b_2/decoder_0/AND_2/B ALU_1b_2/AND_12/w_64_45# 0.06fF
C1868 vdd ALU_1b_2/NOR_2/A 0.03fF
C1869 gnd ALU_1b_2/comparator_0/AND_5/B 0.07fF
C1870 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_6/out 0.05fF
C1871 ALU_1b_3/AND_9/A B2 0.28fF
C1872 vdd ALU_1b_1/AND_2/B 0.10fF
C1873 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.01fF
C1874 ALU_1b_1/AND_0/out ALU_1b_1/AND_2/a_78_51# 0.10fF
C1875 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/A 0.13fF
C1876 ALU_1b_0/AND_7/out gnd 0.07fF
C1877 vdd ALU_1b_3/AND_5/w_64_45# 0.15fF
C1878 ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C1879 ALU_1b_3/NOR_4/A gnd 0.23fF
C1880 ALU_1b_0/AND_16/A ALU_1b_0/AND_16/a_78_51# 0.03fF
C1881 vdd ALU_1b_2/decoder_0/AND_1/a_78_51# 0.06fF
C1882 gnd ALU_1b_3/AND_5/a_78_51# 0.07fF
C1883 ALU_1b_3/comparator_0/w_n220_n67# ALU_1b_3/comparator_0/NOR_2/A 0.06fF
C1884 ALU_1b_0/NOT_4/in F0 0.03fF
C1885 gnd ALU_1b_2/AND_9/a_78_51# 0.07fF
C1886 A2 ALU_1b_3/AND_12/a_78_51# 0.19fF
C1887 ALU_1b_2/AND_0/a_78_51# ALU_1b_2/AND_0/out 0.05fF
C1888 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C1889 ALU_1b_2/AND_1/a_78_51# ALU_1b_2/AND_2/B 0.19fF
C1890 ALU_1b_0/AND_3/out C1 0.01fF
C1891 ALU_1b_2/AND_19/w_64_45# ALU_1b_2/NOR_0/A 0.03fF
C1892 ALU_1b_0/AND_7/w_64_45# ALU_1b_0/AND_7/out 0.03fF
C1893 ALU_1b_0/AND_3/w_64_45# ALU_1b_0/AND_5/B 0.06fF
C1894 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C1895 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.05fF
C1896 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/AND_1/out 0.04fF
C1897 gnd ALU_1b_3/decoder_0/AND_2/B 0.07fF
C1898 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/AND_3/out 0.00fF
C1899 ALU_1b_1/comparator_0/NOR_3/A vdd 0.03fF
C1900 vdd ALU_1b_3/NOR_4/w_n27_1# 0.24fF
C1901 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.03fF
C1902 ALU_1b_1/AND_8/w_64_45# ALU_1b_1/AND_8/a_78_51# 0.09fF
C1903 ALU_1b_2/AND_0/out ALU_1b_2/AND_2/B 0.11fF
C1904 ALU_1b_1/AND_11/a_78_51# ALU_1b_1/AND_9/A 0.03fF
C1905 ALU_1b_1/AND_9/A ALU_1b_1/AND_11/B 0.37fF
C1906 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# vdd 0.14fF
C1907 ALU_1b_3/NOT_2/in ALU_1b_3/NOR_2/A 0.03fF
C1908 ALU_1b_0/NOT_6/in ALU_1b_0/NOR_1/A 0.37fF
C1909 ALU_1b_1/AND_1/out ALU_1b_1/C0 0.01fF
C1910 vdd ALU_1b_3/comparator_0/AND_0/w_64_45# 0.14fF
C1911 ALU_1b_2/comparator_0/AND_3/w_64_45# ALU_1b_2/comparator_0/AND_3/a_78_51# 0.09fF
C1912 ALU_1b_2/AND_9/out ALU_1b_2/AND_7/out 0.02fF
C1913 ALU_1b_2/AND_12/a_78_51# ALU_1b_2/AND_15/A 0.05fF
C1914 ALU_1b_1/AND_12/w_64_45# ALU_1b_1/decoder_0/AND_1/B 0.03fF
C1915 gnd ALU_1b_3/NOT_3/in 0.07fF
C1916 ALU_1b_3/NOT_1/in ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.13fF
C1917 ALU_1b_3/NOR_0/A ALU_1b_3/NOR_3/A 0.01fF
C1918 ALU_1b_0/AND_14/B ALU_1b_0/AND_12/w_64_45# 0.03fF
C1919 gnd ALU_1b_3/comparator_0/AND_0/a_78_51# 0.07fF
C1920 S1 ALU_1b_3/decoder_0/AND_1/B 0.29fF
C1921 ALU_1b_1/comparator_0/AND_3/w_64_45# ALU_1b_1/AND_8/out 0.16fF
C1922 ALU_1b_3/AND_7/a_78_51# ALU_1b_3/AND_8/out 0.10fF
C1923 ALU_1b_0/AND_4/a_78_51# B0 0.03fF
C1924 ALU_1b_3/AND_9/a_78_51# ALU_1b_3/AND_9/out 0.05fF
C1925 ALU_1b_1/NOT_6/in ALU_1b_1/NOR_4/w_n27_1# 0.11fF
C1926 ALU_1b_3/comparator_0/w_113_n67# ALU_1b_3/AND_10/B 0.03fF
C1927 ALU_1b_1/AND_7/a_78_51# vdd 0.06fF
C1928 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/AND_1/out 0.70fF
C1929 ALU_1b_0/AND_5/out gnd 0.62fF
C1930 ALU_1b_0/AND_19/a_78_51# vdd 0.06fF
C1931 gnd ALU_1b_2/C0 0.65fF
C1932 ALU_1b_3/AND_4/w_64_45# B2 0.10fF
C1933 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# vdd 0.06fF
C1934 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out gnd 0.04fF
C1935 ALU_1b_0/comparator_0/AND_4/w_64_45# ALU_1b_0/AND_7/out 0.10fF
C1936 ALU_1b_0/AND_14/A ALU_1b_0/AND_15/A 0.10fF
C1937 ALU_1b_2/comparator_0/NOR_0/A ALU_1b_2/comparator_0/NOR_0/out 0.03fF
C1938 ALU_1b_1/full_adder_1/NOR_0/out ALU_1b_1/AND_18/A 0.04fF
C1939 ALU_1b_0/AND_16/A gnd 0.14fF
C1940 ALU_1b_2/full_adder_0/half_adder_0/w_36_45# ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.09fF
C1941 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.00fF
C1942 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/w_n39_45# 0.11fF
C1943 ALU_1b_2/AND_3/out ALU_1b_2/C0 0.01fF
C1944 ALU_1b_1/AND_14/w_64_45# vdd 0.29fF
C1945 ALU_1b_1/AND_9/out ALU_1b_1/comparator_0/w_n39_45# 0.15fF
C1946 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# vdd 0.14fF
C1947 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_1/AND_1/out 0.04fF
C1948 ALU_1b_1/AND_13/a_78_51# gnd 0.07fF
C1949 ALU_1b_0/decoder_0/AND_3/a_78_51# S1 0.19fF
C1950 vdd ALU_1b_3/AND_15/A 0.43fF
C1951 ALU_1b_3/AND_4/out ALU_1b_3/AND_5/a_78_51# 0.24fF
C1952 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/w_n74_45# 0.03fF
C1953 ALU_1b_0/AND_8/out ALU_1b_0/AND_9/A 0.12fF
C1954 F0 ALU_1b_2/AND_9/a_78_51# 0.19fF
C1955 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_15/B 0.03fF
C1956 ALU_1b_2/AND_13/a_78_51# ALU_1b_2/AND_14/B 0.10fF
C1957 ALU_1b_1/decoder_0/AND_1/B gnd 0.07fF
C1958 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.06fF
C1959 ALU_1b_3/AND_8/out ALU_1b_3/comparator_0/AND_4/a_78_51# 0.20fF
C1960 ALU_1b_1/comparator_0/AND_4/a_78_51# vdd 0.06fF
C1961 ALU_1b_3/AND_15/B ALU_1b_3/AND_15/A 0.28fF
C1962 ALU_1b_1/AND_14/A ALU_1b_1/AND_14/a_78_51# 0.03fF
C1963 ALU_1b_3/AND_6/w_64_45# ALU_1b_3/decoder_0/AND_2/B 0.09fF
C1964 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.09fF
C1965 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_10/a_78_51# 0.09fF
C1966 ALU_1b_0/comparator_0/w_n220_n67# vdd 0.12fF
C1967 ALU_1b_0/AND_0/out Cin 0.01fF
C1968 ALU_1b_1/AND_3/a_78_51# ALU_1b_1/AND_5/B 0.29fF
C1969 ALU_1b_1/AND_9/A gnd 0.35fF
C1970 vdd ALU_1b_3/decoder_0/AND_2/a_78_51# 0.06fF
C1971 ALU_1b_1/NOT_1/in ALU_1b_1/NOT_1/w_n36_43# 0.06fF
C1972 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.20fF
C1973 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_3/AND_3/out 0.13fF
C1974 ALU_1b_0/AND_15/w_64_45# ALU_1b_0/AND_15/a_78_51# 0.09fF
C1975 ALU_1b_0/full_adder_0/w_448_45# vdd 0.12fF
C1976 ALU_1b_1/AND_16/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.03fF
C1977 ALU_1b_1/comparator_0/w_113_n67# ALU_1b_1/comparator_0/NOR_1/out 0.11fF
C1978 ALU_1b_0/AND_3/out vdd 0.03fF
C1979 ALU_1b_1/AND_18/A vdd 0.02fF
C1980 ALU_1b_2/AND_17/A ALU_1b_2/full_adder_0/w_448_45# 0.03fF
C1981 gnd ALU_1b_2/comparator_0/NOR_3/B 0.21fF
C1982 S1 ALU_1b_1/AND_6/w_64_45# 0.62fF
C1983 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/C0 0.19fF
C1984 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# ALU_1b_1/full_adder_1/NOR_0/B 0.36fF
C1985 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.05fF
C1986 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/NOT_1/in 0.13fF
C1987 ALU_1b_0/AND_6/a_78_51# vdd 0.06fF
C1988 ALU_1b_1/AND_3/a_78_51# gnd 0.07fF
C1989 ALU_1b_0/comparator_0/AND_0/w_64_45# ALU_1b_0/AND_6/out 0.26fF
C1990 ALU_1b_0/AND_9/out gnd 0.07fF
C1991 ALU_1b_1/AND_16/A ALU_1b_1/AND_16/a_78_51# 0.03fF
C1992 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_2/a_n14_7# 0.00fF
C1993 ALU_1b_1/NOR_4/B vdd 0.03fF
C1994 F0 ALU_1b_2/C0 8.21fF
C1995 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/AND_1/out 0.06fF
C1996 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_74# 0.02fF
C1997 gnd ALU_1b_3/NOR_0/B 0.17fF
C1998 ALU_1b_1/AND_19/A vdd 0.03fF
C1999 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C2000 ALU_1b_1/AND_2/out ALU_1b_1/AND_2/w_64_45# 0.03fF
C2001 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_9/out 0.19fF
C2002 gnd ALU_1b_3/AND_1/out 0.69fF
C2003 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/NOR_3/out 0.15fF
C2004 ALU_1b_0/AND_8/w_64_45# vdd 0.14fF
C2005 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_0/out 0.23fF
C2006 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C2007 ALU_1b_3/AND_11/a_78_51# ALU_1b_3/AND_11/B 0.19fF
C2008 ALU_1b_1/AND_4/w_64_45# ALU_1b_1/AND_5/B 0.06fF
C2009 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_36# 0.03fF
C2010 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/NOR_0/A 0.16fF
C2011 ALU_1b_0/NOT_3/in ALU_1b_0/NOR_2/B 0.03fF
C2012 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C2013 ALU_1b_0/AND_8/a_78_51# gnd 0.07fF
C2014 ALU_1b_0/comparator_0/AND_0/a_78_51# ALU_1b_0/comparator_0/NOR_0/A 0.05fF
C2015 A1 ALU_1b_2/AND_6/a_78_51# 0.19fF
C2016 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.00fF
C2017 vdd B2 0.21fF
C2018 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd 0.06fF
C2019 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out 0.09fF
C2020 ALU_1b_1/AND_17/w_64_45# ALU_1b_1/NOR_3/B 0.07fF
C2021 ALU_1b_1/AND_8/out ALU_1b_1/C0 0.01fF
C2022 ALU_1b_2/AND_6/w_64_45# ALU_1b_2/decoder_0/AND_1/B 0.13fF
C2023 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_0/a_78_51# 0.29fF
C2024 ALU_1b_3/comparator_0/AND_0/w_64_45# ALU_1b_3/comparator_0/NOR_0/A 0.03fF
C2025 gnd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.14fF
C2026 ALU_1b_0/full_adder_1/NOR_0/B vdd 0.91fF
C2027 ALU_1b_0/comparator_0/AND_5/a_78_51# vdd 0.06fF
C2028 ALU_1b_2/NOR_2/w_n27_1# F1 0.03fF
C2029 ALU_1b_1/AND_3/A ALU_1b_1/AND_5/B 0.42fF
C2030 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.70fF
C2031 ALU_1b_0/AND_19/A ALU_1b_0/AND_19/a_78_51# 0.03fF
C2032 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# ALU_1b_2/full_adder_1/half_adder_1/A 0.06fF
C2033 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_5/B 0.16fF
C2034 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out 0.05fF
C2035 ALU_1b_2/AND_9/A ALU_1b_2/AND_6/w_64_45# 0.36fF
C2036 ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/AND_2/a_78_51# 0.03fF
C2037 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/comparator_0/AND_5/a_78_51# 0.05fF
C2038 ALU_1b_2/full_adder_1/NOR_0/A gnd 0.07fF
C2039 ALU_1b_2/AND_9/w_64_45# F0 0.06fF
C2040 ALU_1b_0/NOR_1/A gnd 0.51fF
C2041 vdd ALU_1b_2/AND_7/out 0.34fF
C2042 ALU_1b_0/AND_10/a_78_51# ALU_1b_0/NOR_1/A 0.05fF
C2043 ALU_1b_2/AND_16/w_64_45# ALU_1b_2/AND_2/B 0.10fF
C2044 ALU_1b_3/AND_19/w_64_45# ALU_1b_3/AND_19/A 0.06fF
C2045 ALU_1b_2/NOT_1/in ALU_1b_2/AND_18/A 0.12fF
C2046 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C2047 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_74# 0.01fF
C2048 ALU_1b_0/AND_12/a_78_51# ALU_1b_0/AND_12/w_64_45# 0.09fF
C2049 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_5/w_64_45# 0.03fF
C2050 ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/AND_2/w_64_45# 0.16fF
C2051 ALU_1b_1/comparator_0/AND_2/w_64_45# ALU_1b_1/comparator_0/AND_2/a_78_51# 0.09fF
C2052 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_4/w_64_45# 0.03fF
C2053 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/AND_7/out 0.11fF
C2054 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/NOR_1/A 0.03fF
C2055 ALU_1b_3/NOR_2/A ALU_1b_3/NOT_3/in 0.23fF
C2056 ALU_1b_0/AND_2/out gnd 0.07fF
C2057 ALU_1b_2/NOR_0/B ALU_1b_2/NOR_3/A 0.01fF
C2058 ALU_1b_1/AND_3/A gnd 0.07fF
C2059 ALU_1b_0/comparator_0/AND_3/w_64_45# ALU_1b_0/comparator_0/AND_5/B 0.06fF
C2060 ALU_1b_3/AND_0/out B2 0.01fF
C2061 ALU_1b_0/NOR_2/B ALU_1b_0/NOR_2/w_n27_1# 0.09fF
C2062 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_0/NAND_0/a_n7_n34# 0.00fF
C2063 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_74# ALU_1b_1/NOT_1/in 0.03fF
C2064 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/AND_3/out 0.14fF
C2065 ALU_1b_0/AND_2/B S1 0.03fF
C2066 ALU_1b_2/NOT_1/in ALU_1b_2/AND_19/A 0.03fF
C2067 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_2/full_adder_1/half_adder_1/A 0.03fF
C2068 ALU_1b_2/AND_16/A gnd 0.14fF
C2069 ALU_1b_1/NOT_1/in ALU_1b_1/full_adder_1/half_adder_1/A 0.23fF
C2070 ALU_1b_2/NOR_4/A ALU_1b_2/NOT_6/in 0.03fF
C2071 ALU_1b_3/AND_19/a_78_51# ALU_1b_3/NOR_0/A 0.16fF
C2072 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_0/AND_16/A 0.03fF
C2073 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/AND_1/out 0.70fF
C2074 ALU_1b_0/AND_5/a_78_51# Cin 0.03fF
C2075 ALU_1b_3/full_adder_1/half_adder_1/w_36_45# ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out 0.09fF
C2076 ALU_1b_1/AND_7/a_78_51# ALU_1b_1/AND_7/out 0.16fF
C2077 ALU_1b_2/C0 ALU_1b_2/AND_2/B 0.28fF
C2078 gnd ALU_1b_2/NOR_1/B 0.22fF
C2079 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_4/a_78_8# 0.00fF
C2080 ALU_1b_1/comparator_0/NOR_2/out vdd 0.03fF
C2081 S1 ALU_1b_1/decoder_0/AND_1/a_78_51# 0.03fF
C2082 ALU_1b_0/comparator_0/w_n39_45# vdd 0.05fF
C2083 ALU_1b_1/AND_2/out ALU_1b_1/AND_1/out 0.11fF
C2084 ALU_1b_2/full_adder_1/half_adder_0/w_36_45# ALU_1b_2/AND_4/out 0.29fF
C2085 ALU_1b_3/AND_5/w_64_45# ALU_1b_3/C0 0.10fF
C2086 ALU_1b_0/full_adder_0/NOR_0/out vdd 0.03fF
C2087 ALU_1b_3/AND_12/w_64_45# ALU_1b_3/AND_5/B 0.03fF
C2088 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C2089 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.09fF
C2090 ALU_1b_2/AND_9/A ALU_1b_2/AND_10/B 0.29fF
C2091 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_74# 0.03fF
C2092 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out gnd 0.04fF
C2093 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.09fF
C2094 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/full_adder_1/w_448_45# 0.11fF
C2095 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOR_3/B 0.20fF
C2096 ALU_1b_0/AND_16/A ALU_1b_0/AND_1/out 0.11fF
C2097 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_0/NOR_0/A 0.06fF
C2098 S1 vdd 3.29fF
C2099 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/w_n74_45# 0.18fF
C2100 ALU_1b_1/AND_12/a_78_51# ALU_1b_1/AND_14/B 0.05fF
C2101 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.05fF
C2102 ALU_1b_3/AND_3/a_78_51# ALU_1b_3/AND_3/A 0.03fF
C2103 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.10fF
C2104 ALU_1b_3/NOR_2/A ALU_1b_3/NOR_2/w_n27_1# 0.06fF
C2105 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C2106 ALU_1b_2/comparator_0/AND_3/a_78_51# ALU_1b_2/AND_8/out 0.03fF
C2107 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/comparator_0/AND_4/a_78_51# 0.04fF
C2108 ALU_1b_2/AND_1/w_64_45# ALU_1b_2/AND_1/out 0.03fF
C2109 ALU_1b_0/comparator_0/NOR_1/A ALU_1b_0/comparator_0/NOR_1/B 0.33fF
C2110 ALU_1b_0/AND_13/a_78_51# ALU_1b_0/AND_14/A 0.05fF
C2111 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/half_adder_1/A 0.01fF
C2112 gnd ALU_1b_3/comparator_0/NOR_1/A 0.17fF
C2113 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/full_adder_1/NOR_0/B 0.05fF
C2114 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# 0.05fF
C2115 ALU_1b_0/AND_4/w_64_45# ALU_1b_0/AND_4/a_78_51# 0.09fF
C2116 ALU_1b_2/decoder_0/AND_1/a_78_51# ALU_1b_2/decoder_0/AND_1/B 0.19fF
C2117 ALU_1b_1/AND_2/out ALU_1b_1/C0 0.16fF
C2118 ALU_1b_2/AND_5/out gnd 0.62fF
C2119 ALU_1b_1/AND_7/out ALU_1b_1/comparator_0/AND_4/a_78_51# 0.03fF
C2120 ALU_1b_3/AND_14/w_64_45# ALU_1b_3/AND_14/A 0.09fF
C2121 ALU_1b_2/AND_4/out ALU_1b_2/AND_4/w_64_45# 0.03fF
C2122 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_2/AND_3/out 0.03fF
C2123 ALU_1b_2/full_adder_0/half_adder_0/w_36_45# vdd 0.14fF
C2124 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_74# vdd 0.02fF
C2125 ALU_1b_1/AND_3/out ALU_1b_1/AND_5/w_64_45# 0.20fF
C2126 ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/AND_2/B 0.05fF
C2127 ALU_1b_1/full_adder_0/NOR_0/B vdd 0.91fF
C2128 ALU_1b_2/NOT_5/in ALU_1b_2/NOR_4/w_n27_1# 0.11fF
C2129 vdd ALU_1b_3/AND_13/a_78_51# 0.06fF
C2130 ALU_1b_2/decoder_0/AND_1/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C2131 ALU_1b_2/AND_3/out ALU_1b_2/AND_5/out 0.11fF
C2132 ALU_1b_0/AND_12/w_64_45# S0 0.68fF
C2133 vdd ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.06fF
C2134 gnd ALU_1b_3/AND_8/out 0.23fF
C2135 vdd ALU_1b_3/decoder_0/AND_1/B 0.03fF
C2136 ALU_1b_1/comparator_0/NOR_0/B ALU_1b_1/comparator_0/w_113_n67# 0.02fF
C2137 ALU_1b_1/comparator_0/w_88_n67# ALU_1b_1/comparator_0/NOR_1/B 0.19fF
C2138 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# 0.04fF
C2139 ALU_1b_1/AND_14/B vdd 0.03fF
C2140 ALU_1b_0/AND_5/out C0 0.01fF
C2141 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/full_adder_1/NOR_0/B 0.00fF
C2142 ALU_1b_0/full_adder_0/NOR_0/A ALU_1b_0/full_adder_0/w_448_45# 0.06fF
C2143 ALU_1b_1/comparator_0/NOR_1/B gnd 0.07fF
C2144 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_2/AND_1/out 0.10fF
C2145 vdd ALU_1b_3/AND_15/w_64_45# 0.15fF
C2146 ALU_1b_1/AND_15/B gnd 0.27fF
C2147 ALU_1b_1/decoder_0/AND_0/a_78_51# ALU_1b_1/decoder_0/AND_2/B 0.03fF
C2148 vdd ALU_1b_3/AND_9/A 1.07fF
C2149 F0 ALU_1b_2/NOR_1/B 0.01fF
C2150 ALU_1b_0/AND_5/B S0 0.03fF
C2151 ALU_1b_0/AND_15/B ALU_1b_0/AND_15/a_78_51# 0.19fF
C2152 ALU_1b_0/AND_2/out ALU_1b_0/AND_2/w_64_45# 0.03fF
C2153 ALU_1b_2/AND_19/w_64_45# ALU_1b_2/AND_5/B 0.06fF
C2154 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.06fF
C2155 ALU_1b_0/comparator_0/w_n220_n67# ALU_1b_0/comparator_0/NOR_2/out 0.11fF
C2156 gnd ALU_1b_3/AND_15/a_78_51# 0.07fF
C2157 ALU_1b_3/AND_7/out ALU_1b_3/comparator_0/w_n74_45# 0.10fF
C2158 ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/NOR_0/out 0.15fF
C2159 ALU_1b_1/AND_1/a_78_51# gnd 0.07fF
C2160 ALU_1b_3/AND_15/B ALU_1b_3/AND_15/w_64_45# 0.06fF
C2161 ALU_1b_3/NOR_1/B ALU_1b_3/NOR_1/A 0.33fF
C2162 ALU_1b_0/NOR_4/A vdd 0.10fF
C2163 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/AND_3/out 0.13fF
C2164 ALU_1b_3/comparator_0/w_n220_n67# ALU_1b_3/comparator_0/NOR_2/B 0.62fF
C2165 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out vdd 0.06fF
C2166 gnd A1 0.48fF
C2167 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.06fF
C2168 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/AND_0/out 0.10fF
C2169 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_2/AND_1/out 0.00fF
C2170 ALU_1b_0/AND_2/out ALU_1b_0/AND_2/a_78_51# 0.05fF
C2171 ALU_1b_0/decoder_0/AND_3/a_78_51# vdd 0.06fF
C2172 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C2173 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/NOR_0/out 0.15fF
C2174 ALU_1b_0/AND_16/w_64_45# ALU_1b_0/NOR_0/B 0.03fF
C2175 vdd ALU_1b_3/AND_3/a_78_51# 0.06fF
C2176 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C2177 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/full_adder_1/half_adder_1/A 0.13fF
C2178 ALU_1b_0/AND_4/out ALU_1b_0/AND_4/w_64_45# 0.03fF
C2179 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/NOR_3/B 0.43fF
C2180 ALU_1b_1/AND_0/out gnd 0.11fF
C2181 ALU_1b_2/AND_7/out B1 0.28fF
C2182 vdd ALU_1b_2/AND_9/out 0.86fF
C2183 S1 ALU_1b_2/decoder_0/AND_2/a_78_51# 0.02fF
C2184 ALU_1b_1/full_adder_0/NOR_0/out gnd 0.07fF
C2185 vdd ALU_1b_3/full_adder_1/half_adder_0/w_36_45# 0.14fF
C2186 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOT_6/in 0.11fF
C2187 C1 ALU_1b_0/AND_2/B 0.01fF
C2188 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C2189 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C2190 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C2191 ALU_1b_0/AND_3/out ALU_1b_0/AND_3/w_64_45# 0.09fF
C2192 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_0/a_78_51# 0.14fF
C2193 gnd ALU_1b_2/NOT_2/in 0.07fF
C2194 ALU_1b_1/decoder_0/AND_1/a_78_51# ALU_1b_1/AND_6/w_64_45# 0.09fF
C2195 ALU_1b_0/NOR_0/w_n27_1# vdd 0.12fF
C2196 ALU_1b_2/AND_5/out F0 0.01fF
C2197 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/full_adder_0/NOR_0/B 0.00fF
C2198 ALU_1b_0/AND_0/a_78_51# A0 0.19fF
C2199 ALU_1b_2/comparator_0/AND_0/w_64_45# ALU_1b_2/AND_9/out 0.30fF
C2200 ALU_1b_0/comparator_0/AND_1/w_64_45# ALU_1b_0/comparator_0/AND_1/a_78_51# 0.09fF
C2201 gnd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# 0.02fF
C2202 ALU_1b_0/AND_15/A gnd 0.87fF
C2203 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C2204 vdd ALU_1b_2/AND_8/a_78_51# 0.06fF
C2205 ALU_1b_2/AND_4/a_78_51# ALU_1b_2/AND_5/B 0.29fF
C2206 ALU_1b_3/full_adder_0/half_adder_1/w_36_45# ALU_1b_3/AND_1/out 0.29fF
C2207 ALU_1b_3/AND_8/out ALU_1b_3/AND_6/w_64_45# 0.15fF
C2208 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# ALU_1b_1/AND_16/A 0.03fF
C2209 ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/decoder_0/AND_1/B 0.29fF
C2210 vdd ALU_1b_1/AND_6/w_64_45# 0.48fF
C2211 ALU_1b_1/decoder_0/AND_3/a_78_51# S0 0.03fF
C2212 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_4/out 0.10fF
C2213 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_1/NOR_0/B 0.52fF
C2214 C1 vdd 0.25fF
C2215 ALU_1b_1/AND_4/out vdd 0.35fF
C2216 ALU_1b_2/AND_17/a_78_51# ALU_1b_2/NOR_3/B 0.07fF
C2217 ALU_1b_0/AND_1/out ALU_1b_0/AND_2/out 0.11fF
C2218 ALU_1b_2/AND_16/A ALU_1b_2/AND_2/B 0.26fF
C2219 ALU_1b_0/decoder_0/AND_2/a_78_51# gnd 0.07fF
C2220 vdd ALU_1b_3/AND_4/w_64_45# 0.15fF
C2221 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_2/A 0.33fF
C2222 vdd ALU_1b_2/NOR_1/A 0.22fF
C2223 ALU_1b_0/AND_0/a_78_51# ALU_1b_0/AND_0/out 0.05fF
C2224 gnd ALU_1b_3/AND_4/a_78_51# 0.07fF
C2225 ALU_1b_3/NOT_4/in ALU_1b_3/NOR_2/w_n27_1# 0.11fF
C2226 gnd ALU_1b_2/AND_14/a_78_51# 0.07fF
C2227 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_4/B 0.03fF
C2228 ALU_1b_1/decoder_0/AND_3/a_78_51# ALU_1b_1/AND_15/A 0.05fF
C2229 ALU_1b_2/NOR_4/w_n27_1# ALU_1b_2/NOR_1/A 0.09fF
C2230 ALU_1b_0/comparator_0/NOR_0/out vdd 0.03fF
C2231 ALU_1b_2/AND_3/w_64_45# A1 0.10fF
C2232 ALU_1b_3/AND_16/a_78_51# ALU_1b_3/AND_2/B 0.19fF
C2233 ALU_1b_3/full_adder_1/NOR_0/B gnd 0.07fF
C2234 ALU_1b_3/C0 B2 2.32fF
C2235 vdd ALU_1b_3/AND_3/A 0.03fF
C2236 ALU_1b_2/comparator_0/NOR_3/B ALU_1b_2/comparator_0/AND_4/a_78_51# 0.18fF
C2237 ALU_1b_2/NOT_2/in ALU_1b_2/NOR_0/w_n27_1# 0.11fF
C2238 ALU_1b_0/AND_6/out ALU_1b_0/AND_9/A 0.01fF
C2239 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_74# vdd 0.02fF
C2240 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.09fF
C2241 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_1/AND_5/out 0.05fF
C2242 C0 ALU_1b_0/AND_8/a_78_51# 0.19fF
C2243 ALU_1b_3/AND_18/w_64_45# ALU_1b_3/AND_18/a_78_51# 0.09fF
C2244 ALU_1b_3/NOT_6/in ALU_1b_1/C0 0.03fF
C2245 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/AND_1/out 0.20fF
C2246 ALU_1b_0/full_adder_0/NOR_0/out ALU_1b_0/full_adder_0/NOR_0/A 0.03fF
C2247 ALU_1b_1/comparator_0/AND_3/w_64_45# ALU_1b_1/comparator_0/NOR_2/A 0.03fF
C2248 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_3/a_78_51# 0.19fF
C2249 ALU_1b_1/comparator_0/NOR_0/A ALU_1b_1/comparator_0/w_88_n67# 0.06fF
C2250 ALU_1b_1/comparator_0/AND_2/B vdd 0.03fF
C2251 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C2252 vdd ALU_1b_1/AND_10/B 1.59fF
C2253 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/A 0.06fF
C2254 ALU_1b_3/AND_5/out ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C2255 ALU_1b_1/NOR_2/B gnd 0.07fF
C2256 vdd ALU_1b_3/comparator_0/AND_1/w_64_45# 0.14fF
C2257 ALU_1b_1/comparator_0/NOR_0/A gnd 0.17fF
C2258 ALU_1b_1/full_adder_1/NOR_0/out vdd 0.03fF
C2259 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/AND_8/out 0.38fF
C2260 ALU_1b_0/NOR_1/B ALU_1b_0/NOT_3/in 0.15fF
C2261 ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C2262 ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/AND_10/B 0.09fF
C2263 gnd ALU_1b_3/comparator_0/AND_1/a_78_51# 0.07fF
C2264 B0 gnd 0.38fF
C2265 ALU_1b_3/AND_5/out ALU_1b_3/AND_5/w_64_45# 0.03fF
C2266 ALU_1b_1/comparator_0/AND_5/w_64_45# ALU_1b_1/AND_8/out 0.32fF
C2267 ALU_1b_1/AND_12/a_78_51# vdd 0.06fF
C2268 ALU_1b_1/AND_8/w_64_45# ALU_1b_1/AND_9/A 0.39fF
C2269 F2 ALU_1b_3/NOR_2/w_n27_1# 0.03fF
C2270 ALU_1b_0/AND_18/a_78_51# vdd 0.06fF
C2271 vdd ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C2272 ALU_1b_0/AND_2/out C0 0.01fF
C2273 vdd ALU_1b_1/NOR_2/A 0.03fF
C2274 ALU_1b_1/comparator_0/AND_5/B gnd 0.07fF
C2275 ALU_1b_1/AND_9/A F2 0.28fF
C2276 ALU_1b_1/AND_3/out B3 0.01fF
C2277 ALU_1b_0/AND_2/B vdd 0.10fF
C2278 ALU_1b_0/AND_0/out ALU_1b_0/full_adder_0/NOR_0/B 0.10fF
C2279 vdd ALU_1b_2/AND_5/w_64_45# 0.15fF
C2280 ALU_1b_0/AND_7/w_64_45# B0 0.06fF
C2281 ALU_1b_2/NOR_4/A gnd 0.23fF
C2282 ALU_1b_3/AND_3/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.26fF
C2283 ALU_1b_2/AND_0/a_78_51# A1 0.19fF
C2284 ALU_1b_1/comparator_0/NOR_1/A ALU_1b_1/comparator_0/NOR_1/out 0.03fF
C2285 ALU_1b_1/decoder_0/AND_1/a_78_51# vdd 0.06fF
C2286 gnd ALU_1b_2/AND_5/a_78_51# 0.07fF
C2287 ALU_1b_1/AND_9/a_78_51# gnd 0.07fF
C2288 ALU_1b_2/AND_7/out ALU_1b_2/AND_9/A 0.01fF
C2289 ALU_1b_3/AND_4/out ALU_1b_3/AND_4/a_78_51# 0.05fF
C2290 ALU_1b_0/NOR_1/B ALU_1b_0/NOR_2/w_n27_1# 0.06fF
C2291 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_1/full_adder_1/half_adder_1/A 0.26fF
C2292 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.52fF
C2293 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_6/w_64_45# 0.09fF
C2294 gnd ALU_1b_3/AND_14/A 0.07fF
C2295 A1 ALU_1b_2/AND_2/B 0.50fF
C2296 ALU_1b_2/AND_3/out ALU_1b_2/AND_5/a_78_51# 0.10fF
C2297 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/AND_4/out 0.09fF
C2298 ALU_1b_3/AND_14/A ALU_1b_3/AND_14/B 0.42fF
C2299 ALU_1b_3/AND_9/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C2300 ALU_1b_1/NOR_0/A ALU_1b_1/NOT_2/in 0.03fF
C2301 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/w_448_45# 0.16fF
C2302 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/NOR_0/B 0.48fF
C2303 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_11/a_78_51# 0.09fF
C2304 gnd ALU_1b_2/decoder_0/AND_2/B 0.07fF
C2305 ALU_1b_0/comparator_0/NOR_3/A vdd 0.03fF
C2306 vdd ALU_1b_3/comparator_0/NOR_1/B 0.30fF
C2307 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_11/B 0.11fF
C2308 vdd ALU_1b_2/NOR_4/w_n27_1# 0.24fF
C2309 ALU_1b_2/NOT_1/in ALU_1b_2/full_adder_1/NOR_0/out 0.10fF
C2310 ALU_1b_0/comparator_0/NOR_1/B ALU_1b_0/comparator_0/NOR_1/out 0.25fF
C2311 vdd ALU_1b_3/AND_15/B 0.09fF
C2312 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOT_5/in 0.11fF
C2313 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_16/A 0.23fF
C2314 ALU_1b_0/comparator_0/w_n195_n67# ALU_1b_0/comparator_0/NOR_3/B 0.06fF
C2315 gnd ALU_1b_3/comparator_0/NOR_1/out 0.07fF
C2316 vdd ALU_1b_2/comparator_0/AND_0/w_64_45# 0.14fF
C2317 ALU_1b_1/NOR_4/B ALU_1b_1/NOR_1/A 0.07fF
C2318 ALU_1b_2/AND_17/A ALU_1b_2/AND_17/w_64_45# 0.06fF
C2319 ALU_1b_3/NOR_0/A ALU_1b_3/NOR_0/w_n27_1# 0.06fF
C2320 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C2321 vdd ALU_1b_3/AND_1/a_78_51# 0.06fF
C2322 gnd ALU_1b_2/NOT_3/in 0.07fF
C2323 ALU_1b_3/AND_19/a_78_51# ALU_1b_3/AND_5/B 0.19fF
C2324 gnd ALU_1b_2/comparator_0/AND_0/a_78_51# 0.07fF
C2325 S1 ALU_1b_2/decoder_0/AND_1/B 0.29fF
C2326 ALU_1b_3/comparator_0/w_n220_n67# ALU_1b_3/AND_11/B 0.03fF
C2327 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out ALU_1b_1/AND_5/out 0.08fF
C2328 ALU_1b_0/AND_7/a_78_51# vdd 0.06fF
C2329 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# ALU_1b_0/AND_2/out 0.29fF
C2330 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# ALU_1b_0/full_adder_0/NOR_0/B 0.36fF
C2331 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_1/w_64_45# 0.10fF
C2332 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/comparator_0/NOR_3/out 0.05fF
C2333 gnd ALU_1b_3/NOR_3/B 0.23fF
C2334 vdd ALU_1b_3/AND_0/out 0.03fF
C2335 vdd ALU_1b_3/full_adder_0/NOR_0/out 0.03fF
C2336 ALU_1b_1/AND_16/a_78_51# ALU_1b_1/NOR_0/B 0.05fF
C2337 vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C2338 ALU_1b_1/AND_7/out ALU_1b_1/AND_6/w_64_45# 0.13fF
C2339 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/NOR_0/out 0.15fF
C2340 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/NOR_3/out 0.03fF
C2341 ALU_1b_3/AND_9/A ALU_1b_3/C0 0.28fF
C2342 ALU_1b_0/AND_2/w_64_45# B0 0.10fF
C2343 ALU_1b_0/AND_14/w_64_45# vdd 0.29fF
C2344 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/full_adder_1/NOR_0/A 0.05fF
C2345 ALU_1b_2/AND_0/w_64_45# ALU_1b_2/AND_0/a_78_51# 0.09fF
C2346 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/NOR_0/out 0.03fF
C2347 ALU_1b_3/full_adder_1/w_448_45# ALU_1b_3/AND_18/A 0.03fF
C2348 ALU_1b_1/NOR_2/A ALU_1b_1/NOT_4/in 0.03fF
C2349 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out 0.05fF
C2350 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_2/full_adder_1/half_adder_1/A 0.03fF
C2351 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C2352 ALU_1b_3/AND_2/out F1 0.01fF
C2353 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.52fF
C2354 ALU_1b_0/AND_18/A ALU_1b_0/AND_18/a_78_51# 0.03fF
C2355 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out 0.05fF
C2356 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/NOR_0/A 0.12fF
C2357 ALU_1b_0/AND_13/a_78_51# gnd 0.07fF
C2358 vdd ALU_1b_2/AND_15/A 0.43fF
C2359 ALU_1b_3/AND_0/out ALU_1b_3/AND_1/a_78_51# 0.10fF
C2360 ALU_1b_3/NOR_4/A ALU_1b_3/NOR_1/A 0.01fF
C2361 ALU_1b_3/AND_18/A ALU_1b_3/AND_18/w_64_45# 0.06fF
C2362 ALU_1b_0/AND_2/a_78_51# B0 0.03fF
C2363 ALU_1b_0/decoder_0/AND_1/B gnd 0.07fF
C2364 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_1/a_78_51# 0.10fF
C2365 ALU_1b_3/comparator_0/AND_0/a_78_51# ALU_1b_3/AND_9/out 0.02fF
C2366 ALU_1b_3/AND_7/w_64_45# ALU_1b_3/AND_7/a_78_51# 0.09fF
C2367 ALU_1b_0/comparator_0/AND_4/a_78_51# vdd 0.06fF
C2368 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_1/AND_4/out 0.06fF
C2369 ALU_1b_2/AND_0/w_64_45# ALU_1b_2/AND_2/B 0.06fF
C2370 ALU_1b_3/NOR_1/B B2 0.01fF
C2371 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.70fF
C2372 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/NOR_0/B 0.00fF
C2373 ALU_1b_2/AND_19/w_64_45# ALU_1b_2/AND_19/a_78_51# 0.09fF
C2374 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out vdd 0.06fF
C2375 ALU_1b_0/comparator_0/AND_2/w_64_45# ALU_1b_0/comparator_0/NOR_1/A 0.03fF
C2376 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/AND_8/out 0.02fF
C2377 ALU_1b_0/AND_9/A gnd 0.35fF
C2378 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/AND_3/out 0.14fF
C2379 vdd ALU_1b_2/decoder_0/AND_2/a_78_51# 0.06fF
C2380 ALU_1b_0/AND_10/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C2381 ALU_1b_2/AND_17/w_64_45# ALU_1b_2/AND_2/B 0.06fF
C2382 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.01fF
C2383 ALU_1b_2/NOR_2/A ALU_1b_2/NOR_2/B 0.47fF
C2384 ALU_1b_0/NOR_1/A ALU_1b_0/AND_11/B 0.03fF
C2385 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_1/full_adder_1/half_adder_1/A 0.03fF
C2386 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# ALU_1b_1/AND_2/out 0.29fF
C2387 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/AND_16/A 0.06fF
C2388 gnd ALU_1b_3/decoder_0/AND_0/a_78_51# 0.07fF
C2389 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# gnd 0.11fF
C2390 ALU_1b_1/AND_6/out ALU_1b_1/AND_8/out 0.10fF
C2391 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/AND_7/out 0.05fF
C2392 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C2393 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_9/A 0.95fF
C2394 A2 ALU_1b_3/AND_15/A 0.42fF
C2395 ALU_1b_2/AND_2/out ALU_1b_2/AND_2/a_78_51# 0.05fF
C2396 ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/comparator_0/NOR_2/A 0.03fF
C2397 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_2/NOT_1/in 0.03fF
C2398 ALU_1b_0/AND_18/A vdd 0.02fF
C2399 ALU_1b_1/AND_5/out ALU_1b_1/full_adder_1/half_adder_1/A 0.72fF
C2400 ALU_1b_3/AND_2/a_78_51# ALU_1b_3/AND_2/B 0.29fF
C2401 ALU_1b_2/NOR_3/B ALU_1b_2/NOR_3/A 0.34fF
C2402 ALU_1b_0/AND_6/w_64_45# S1 0.62fF
C2403 ALU_1b_1/comparator_0/NOR_3/B gnd 0.21fF
C2404 ALU_1b_0/comparator_0/AND_1/w_64_45# ALU_1b_0/comparator_0/NOR_0/B 0.03fF
C2405 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_5/w_64_45# 0.06fF
C2406 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_8/out 0.11fF
C2407 ALU_1b_0/AND_7/w_64_45# ALU_1b_0/AND_9/A 0.39fF
C2408 B3 ALU_1b_1/AND_2/B 0.28fF
C2409 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_74# vdd 0.02fF
C2410 ALU_1b_0/AND_3/a_78_51# gnd 0.07fF
C2411 gnd ALU_1b_3/AND_6/out 0.07fF
C2412 ALU_1b_3/NOR_1/A ALU_1b_3/NOT_3/in 0.03fF
C2413 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.01fF
C2414 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_4/a_78_8# 0.00fF
C2415 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_15/A 0.50fF
C2416 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_74# vdd 0.02fF
C2417 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C2418 gnd ALU_1b_2/NOR_0/B 0.17fF
C2419 ALU_1b_2/AND_4/out ALU_1b_2/C0 0.16fF
C2420 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_3/NOT_1/in 0.03fF
C2421 ALU_1b_0/AND_19/A vdd 0.03fF
C2422 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.08fF
C2423 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_1/NOT_1/in 0.03fF
C2424 ALU_1b_1/AND_3/out ALU_1b_1/AND_3/a_78_51# 0.05fF
C2425 vdd ALU_1b_3/NOR_2/B 0.03fF
C2426 S0 ALU_1b_3/decoder_0/AND_2/a_78_51# 0.05fF
C2427 ALU_1b_1/NOR_4/B ALU_1b_1/NOR_4/w_n27_1# 0.09fF
C2428 ALU_1b_2/AND_1/out gnd 0.69fF
C2429 ALU_1b_2/AND_8/w_64_45# ALU_1b_2/AND_8/out 0.03fF
C2430 vdd ALU_1b_3/comparator_0/NOR_0/A 0.03fF
C2431 ALU_1b_2/comparator_0/AND_3/a_78_51# ALU_1b_2/comparator_0/NOR_2/A 0.17fF
C2432 ALU_1b_2/AND_9/out ALU_1b_2/AND_9/A 0.04fF
C2433 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C2434 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/comparator_0/w_n39_45# 0.03fF
C2435 ALU_1b_1/full_adder_1/half_adder_0/w_36_45# ALU_1b_1/AND_3/out 0.09fF
C2436 ALU_1b_3/AND_2/out ALU_1b_3/AND_2/B 0.38fF
C2437 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/AND_5/out 0.20fF
C2438 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_74# 0.01fF
C2439 F3 vdd 0.12fF
C2440 vdd B1 0.28fF
C2441 ALU_1b_3/comparator_0/NOR_1/out ALU_1b_3/AND_10/B 0.05fF
C2442 ALU_1b_3/AND_5/w_64_45# ALU_1b_3/AND_5/a_78_51# 0.09fF
C2443 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C2444 vdd ALU_1b_3/comparator_0/AND_5/B 0.03fF
C2445 ALU_1b_2/comparator_0/AND_5/a_78_51# ALU_1b_2/AND_8/out 0.02fF
C2446 ALU_1b_0/AND_1/a_78_51# gnd 0.07fF
C2447 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_14/a_78_51# 0.09fF
C2448 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C2449 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/NOR_0/out 0.03fF
C2450 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_3/AND_4/out 0.70fF
C2451 ALU_1b_0/NOR_0/B ALU_1b_0/NOT_2/in 0.15fF
C2452 ALU_1b_3/AND_3/out ALU_1b_3/full_adder_1/half_adder_1/A 0.23fF
C2453 gnd ALU_1b_3/comparator_0/NOR_2/A 0.24fF
C2454 ALU_1b_3/AND_7/out ALU_1b_3/AND_8/out 0.40fF
C2455 ALU_1b_3/comparator_0/AND_4/w_64_45# ALU_1b_3/comparator_0/AND_4/a_78_51# 0.09fF
C2456 ALU_1b_1/AND_7/out vdd 0.34fF
C2457 ALU_1b_3/AND_14/a_78_51# ALU_1b_3/AND_15/A 0.00fF
C2458 ALU_1b_3/NOR_1/A ALU_1b_3/NOR_2/w_n27_1# 0.10fF
C2459 ALU_1b_3/AND_6/w_64_45# ALU_1b_3/decoder_0/AND_0/a_78_51# 0.09fF
C2460 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_1/half_adder_1/A 0.13fF
C2461 A2 B2 0.64fF
C2462 ALU_1b_1/AND_2/w_64_45# ALU_1b_1/AND_2/a_78_51# 0.09fF
C2463 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.09fF
C2464 ALU_1b_2/comparator_0/w_88_n67# ALU_1b_2/comparator_0/NOR_0/B 0.20fF
C2465 ALU_1b_1/AND_7/a_78_51# B3 0.19fF
C2466 ALU_1b_1/AND_3/out ALU_1b_1/AND_4/w_64_45# 0.20fF
C2467 ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/NOR_1/B 0.01fF
C2468 ALU_1b_2/NOR_0/B ALU_1b_2/NOR_0/w_n27_1# 0.06fF
C2469 ALU_1b_3/NOR_4/A ALU_1b_3/NOR_4/w_n27_1# 0.10fF
C2470 vdd ALU_1b_3/AND_9/a_78_51# 0.06fF
C2471 ALU_1b_2/NOR_1/A ALU_1b_2/AND_9/A 0.03fF
C2472 ALU_1b_0/full_adder_0/NOR_0/A vdd 0.03fF
C2473 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_2/AND_16/A 0.03fF
C2474 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/AND_16/A 0.05fF
C2475 ALU_1b_0/AND_3/A gnd 0.07fF
C2476 ALU_1b_0/AND_4/out Cin 0.15fF
C2477 ALU_1b_1/AND_3/w_64_45# ALU_1b_1/AND_3/a_78_51# 0.09fF
C2478 gnd ALU_1b_3/comparator_0/NOR_0/B 0.17fF
C2479 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# vdd 0.06fF
C2480 ALU_1b_1/AND_0/out F2 0.01fF
C2481 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# vdd 0.22fF
C2482 ALU_1b_1/AND_16/A gnd 0.14fF
C2483 ALU_1b_3/AND_6/out ALU_1b_3/AND_6/w_64_45# 0.14fF
C2484 ALU_1b_1/AND_14/w_64_45# B3 0.06fF
C2485 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/NOT_1/in 0.23fF
C2486 ALU_1b_1/NOR_1/B gnd 0.22fF
C2487 vdd ALU_1b_3/AND_16/w_64_45# 0.15fF
C2488 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C2489 ALU_1b_0/comparator_0/NOR_2/out vdd 0.03fF
C2490 ALU_1b_0/decoder_0/AND_1/a_78_51# S1 0.03fF
C2491 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/w_448_45# 0.16fF
C2492 ALU_1b_0/AND_15/a_78_51# ALU_1b_0/NOR_1/B 0.05fF
C2493 ALU_1b_2/AND_18/w_64_45# ALU_1b_2/AND_5/B 0.10fF
C2494 vdd ALU_1b_3/full_adder_0/w_448_45# 0.12fF
C2495 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_36# gnd 0.02fF
C2496 gnd ALU_1b_3/AND_16/a_78_51# 0.07fF
C2497 ALU_1b_2/AND_15/A B1 0.28fF
C2498 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_10/B 0.20fF
C2499 ALU_1b_2/AND_1/out F0 0.01fF
C2500 ALU_1b_3/AND_15/w_64_45# ALU_1b_3/NOR_1/B 0.06fF
C2501 ALU_1b_0/AND_5/w_64_45# ALU_1b_0/AND_5/B 0.06fF
C2502 ALU_1b_1/full_adder_1/NOR_0/A vdd 0.03fF
C2503 ALU_1b_2/AND_2/w_64_45# ALU_1b_2/AND_2/B 0.06fF
C2504 ALU_1b_0/AND_3/w_64_45# vdd 0.21fF
C2505 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/full_adder_0/w_448_45# 0.06fF
C2506 ALU_1b_1/comparator_0/w_n195_n67# ALU_1b_1/comparator_0/NOR_3/out 0.11fF
C2507 ALU_1b_3/AND_17/A ALU_1b_3/AND_17/a_78_51# 0.03fF
C2508 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_0/AND_5/out 0.10fF
C2509 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C2510 ALU_1b_2/NOT_4/in ALU_1b_2/NOR_2/B 0.15fF
C2511 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# gnd 0.02fF
C2512 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/NOR_0/A 0.10fF
C2513 ALU_1b_1/decoder_0/AND_1/B ALU_1b_1/AND_2/B 0.17fF
C2514 vdd ALU_1b_3/C0 0.44fF
C2515 ALU_1b_1/AND_17/w_64_45# ALU_1b_1/AND_17/a_78_51# 0.09fF
C2516 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.09fF
C2517 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_2/B 0.40fF
C2518 ALU_1b_3/comparator_0/AND_0/w_64_45# ALU_1b_3/comparator_0/AND_0/a_78_51# 0.09fF
C2519 F3 ALU_1b_1/NOT_4/in 0.03fF
C2520 ALU_1b_1/AND_6/out ALU_1b_1/comparator_0/AND_1/a_78_51# 0.03fF
C2521 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/AND_9/out 0.29fF
C2522 ALU_1b_2/NOR_4/w_n27_1# ALU_1b_3/C0 0.03fF
C2523 gnd ALU_1b_2/comparator_0/NOR_1/A 0.17fF
C2524 ALU_1b_0/NOR_4/B ALU_1b_0/NOT_6/in 0.15fF
C2525 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C2526 ALU_1b_1/AND_5/out gnd 0.62fF
C2527 ALU_1b_1/AND_9/out ALU_1b_1/AND_10/B 0.06fF
C2528 A3 ALU_1b_1/AND_12/w_64_45# 0.18fF
C2529 ALU_1b_0/NOT_1/in ALU_1b_0/full_adder_1/NOR_0/A 0.23fF
C2530 ALU_1b_2/comparator_0/AND_1/w_64_45# ALU_1b_2/AND_9/out 0.39fF
C2531 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_2/w_64_45# 0.06fF
C2532 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_5/B 0.05fF
C2533 ALU_1b_3/full_adder_0/w_448_45# ALU_1b_3/full_adder_0/NOR_0/out 0.11fF
C2534 ALU_1b_3/AND_1/a_78_51# ALU_1b_3/C0 0.03fF
C2535 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.04fF
C2536 ALU_1b_1/AND_3/w_64_45# ALU_1b_1/AND_3/A 0.09fF
C2537 vdd ALU_1b_2/AND_13/a_78_51# 0.06fF
C2538 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.03fF
C2539 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.09fF
C2540 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C2541 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out vdd 0.06fF
C2542 ALU_1b_1/NOR_0/B ALU_1b_1/NOR_0/A 0.33fF
C2543 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_1/A 0.11fF
C2544 S1 S0 12.40fF
C2545 gnd ALU_1b_2/AND_8/out 0.23fF
C2546 vdd ALU_1b_2/decoder_0/AND_1/B 0.03fF
C2547 ALU_1b_1/AND_1/w_64_45# ALU_1b_1/AND_2/B 0.06fF
C2548 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C2549 ALU_1b_0/AND_14/B vdd 0.03fF
C2550 ALU_1b_3/decoder_0/AND_3/a_78_51# ALU_1b_3/AND_12/w_64_45# 0.09fF
C2551 A3 ALU_1b_1/AND_5/B 0.01fF
C2552 ALU_1b_3/AND_3/out ALU_1b_3/AND_5/B 0.11fF
C2553 ALU_1b_3/AND_0/out ALU_1b_3/C0 0.01fF
C2554 ALU_1b_0/comparator_0/NOR_1/B gnd 0.07fF
C2555 vdd ALU_1b_3/AND_9/w_64_45# 0.42fF
C2556 ALU_1b_0/NOT_3/in ALU_1b_0/NOR_2/w_n27_1# 0.11fF
C2557 ALU_1b_0/AND_15/B gnd 0.27fF
C2558 A0 ALU_1b_0/AND_8/out 0.11fF
C2559 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_7/out 0.20fF
C2560 vdd ALU_1b_2/AND_15/w_64_45# 0.15fF
C2561 vdd ALU_1b_2/AND_9/A 1.07fF
C2562 ALU_1b_3/AND_19/A ALU_1b_3/NOR_0/A 0.10fF
C2563 ALU_1b_0/AND_15/A ALU_1b_0/AND_12/w_64_45# 0.36fF
C2564 ALU_1b_0/NOR_0/w_n27_1# ALU_1b_0/NOR_2/A 0.03fF
C2565 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_0/AND_16/A 0.13fF
C2566 gnd ALU_1b_3/AND_10/a_78_51# 0.07fF
C2567 ALU_1b_3/decoder_0/AND_2/a_78_51# ALU_1b_3/decoder_0/AND_2/B 0.19fF
C2568 ALU_1b_1/comparator_0/AND_2/a_78_51# ALU_1b_1/comparator_0/NOR_1/A 0.38fF
C2569 gnd ALU_1b_2/AND_15/a_78_51# 0.07fF
C2570 ALU_1b_2/NOR_4/A ALU_1b_2/NOR_4/B 0.35fF
C2571 ALU_1b_3/AND_17/a_78_51# ALU_1b_3/AND_2/B 0.19fF
C2572 ALU_1b_2/AND_18/w_64_45# ALU_1b_2/NOR_3/A 0.03fF
C2573 ALU_1b_2/full_adder_0/half_adder_0/w_36_45# ALU_1b_2/AND_0/out 0.09fF
C2574 A3 gnd 0.48fF
C2575 vdd ALU_1b_3/comparator_0/NOR_3/B 0.03fF
C2576 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/NOR_0/out 0.03fF
C2577 ALU_1b_0/comparator_0/NOR_0/A ALU_1b_0/comparator_0/NOR_0/B 0.33fF
C2578 ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.14fF
C2579 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_74# 0.03fF
C2580 vdd ALU_1b_2/AND_3/a_78_51# 0.06fF
C2581 ALU_1b_0/decoder_0/AND_2/a_78_51# ALU_1b_0/AND_12/w_64_45# 0.09fF
C2582 S0 ALU_1b_3/decoder_0/AND_1/B 0.03fF
C2583 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/NOR_0/B 0.12fF
C2584 gnd ALU_1b_3/comparator_0/NOR_3/out 0.07fF
C2585 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/full_adder_1/NOR_0/A 0.03fF
C2586 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_36# 0.03fF
C2587 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/NOR_0/A 0.16fF
C2588 ALU_1b_0/AND_1/w_64_45# ALU_1b_0/AND_1/out 0.03fF
C2589 ALU_1b_0/AND_6/w_64_45# ALU_1b_0/AND_2/B 0.03fF
C2590 ALU_1b_1/AND_9/out vdd 0.86fF
C2591 ALU_1b_1/comparator_0/AND_1/a_78_51# ALU_1b_1/comparator_0/NOR_0/B 0.05fF
C2592 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_5/a_78_51# 0.29fF
C2593 S1 ALU_1b_1/decoder_0/AND_2/a_78_51# 0.02fF
C2594 A2 ALU_1b_3/AND_9/A 0.31fF
C2595 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_13/a_78_51# 0.09fF
C2596 ALU_1b_1/AND_7/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C2597 ALU_1b_2/full_adder_1/half_adder_0/w_36_45# vdd 0.14fF
C2598 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_74# vdd 0.02fF
C2599 ALU_1b_1/NOR_1/A ALU_1b_1/NOR_2/A 0.12fF
C2600 ALU_1b_1/NOT_2/in gnd 0.07fF
C2601 vdd ALU_1b_3/comparator_0/AND_2/w_64_45# 0.15fF
C2602 ALU_1b_2/comparator_0/AND_5/w_64_45# ALU_1b_2/comparator_0/AND_5/a_78_51# 0.09fF
C2603 ALU_1b_2/comparator_0/AND_5/B ALU_1b_2/AND_7/out 0.61fF
C2604 ALU_1b_0/comparator_0/AND_5/a_78_51# ALU_1b_0/AND_7/out 0.14fF
C2605 ALU_1b_0/comparator_0/NOR_1/A ALU_1b_0/comparator_0/w_113_n67# 0.06fF
C2606 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_14/B 0.06fF
C2607 ALU_1b_1/AND_9/a_78_51# F2 0.19fF
C2608 ALU_1b_2/AND_13/a_78_51# ALU_1b_2/AND_15/A 0.05fF
C2609 C0 ALU_1b_0/AND_9/A 0.28fF
C2610 vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.06fF
C2611 ALU_1b_0/AND_1/out ALU_1b_0/AND_1/a_78_51# 0.05fF
C2612 ALU_1b_2/AND_4/out ALU_1b_2/AND_5/out 0.11fF
C2613 ALU_1b_0/decoder_0/AND_2/a_78_51# ALU_1b_0/AND_5/B 0.05fF
C2614 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/AND_4/out 0.11fF
C2615 ALU_1b_0/AND_5/out ALU_1b_0/AND_3/out 0.11fF
C2616 ALU_1b_3/AND_3/w_64_45# ALU_1b_3/AND_5/B 0.06fF
C2617 ALU_1b_3/comparator_0/AND_5/w_64_45# ALU_1b_3/AND_7/out 0.30fF
C2618 gnd ALU_1b_3/comparator_0/AND_2/a_78_51# 0.07fF
C2619 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C2620 ALU_1b_1/comparator_0/AND_4/w_64_45# ALU_1b_1/AND_8/out 0.37fF
C2621 ALU_1b_3/AND_8/a_78_51# ALU_1b_3/AND_8/out 0.22fF
C2622 ALU_1b_1/AND_8/a_78_51# vdd 0.06fF
C2623 ALU_1b_1/AND_14/B ALU_1b_1/AND_15/A 0.16fF
C2624 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/AND_16/A 0.01fF
C2625 F1 ALU_1b_3/AND_5/B 0.01fF
C2626 ALU_1b_0/AND_6/w_64_45# vdd 0.48fF
C2627 ALU_1b_0/decoder_0/AND_3/a_78_51# S0 0.03fF
C2628 ALU_1b_2/AND_15/w_64_45# ALU_1b_2/AND_15/A 0.06fF
C2629 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# ALU_1b_0/full_adder_1/half_adder_1/A 0.06fF
C2630 vdd ALU_1b_2/AND_4/w_64_45# 0.15fF
C2631 ALU_1b_2/NOR_1/B ALU_1b_2/NOR_2/A 0.00fF
C2632 ALU_1b_3/full_adder_1/w_448_45# ALU_1b_3/full_adder_1/NOR_0/out 0.11fF
C2633 ALU_1b_3/AND_19/A ALU_1b_3/NOT_1/w_n36_43# 0.03fF
C2634 ALU_1b_3/full_adder_1/NOR_0/A vdd 0.03fF
C2635 ALU_1b_1/NOR_1/A vdd 0.22fF
C2636 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_0/NAND_0/a_n7_n34# 0.00fF
C2637 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/AND_0/out 0.14fF
C2638 gnd ALU_1b_2/AND_4/a_78_51# 0.07fF
C2639 ALU_1b_1/AND_14/a_78_51# gnd 0.07fF
C2640 ALU_1b_0/AND_7/out ALU_1b_0/comparator_0/w_n39_45# 0.06fF
C2641 ALU_1b_2/AND_14/B ALU_1b_2/AND_14/a_78_51# 0.19fF
C2642 ALU_1b_2/full_adder_1/NOR_0/B gnd 0.07fF
C2643 A1 ALU_1b_2/AND_6/w_64_45# 0.06fF
C2644 vdd ALU_1b_2/AND_3/A 0.03fF
C2645 ALU_1b_3/comparator_0/w_88_n67# ALU_1b_3/comparator_0/NOR_0/out 0.11fF
C2646 ALU_1b_2/AND_3/out ALU_1b_2/AND_4/a_78_51# 0.10fF
C2647 ALU_1b_1/comparator_0/NOR_0/out ALU_1b_1/comparator_0/NOR_1/B 0.05fF
C2648 ALU_1b_0/AND_5/out ALU_1b_0/full_adder_1/NOR_0/B 0.19fF
C2649 B0 ALU_1b_0/AND_5/B 0.28fF
C2650 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/w_n195_n67# 0.19fF
C2651 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out ALU_1b_0/full_adder_1/NOR_0/B 0.00fF
C2652 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_74# 0.03fF
C2653 ALU_1b_0/comparator_0/AND_2/B vdd 0.03fF
C2654 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/AND_3/out 0.10fF
C2655 ALU_1b_2/comparator_0/NOR_1/B ALU_1b_2/comparator_0/NOR_1/a_n14_7# 0.00fF
C2656 ALU_1b_0/NOR_4/B gnd 0.07fF
C2657 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_2/AND_1/out 0.04fF
C2658 ALU_1b_3/AND_2/w_64_45# B2 0.10fF
C2659 vdd ALU_1b_3/NOR_1/B 0.20fF
C2660 ALU_1b_0/AND_16/w_64_45# ALU_1b_0/AND_16/a_78_51# 0.09fF
C2661 ALU_1b_0/AND_10/B vdd 1.59fF
C2662 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/AND_16/A 0.22fF
C2663 ALU_1b_0/NOR_2/B gnd 0.07fF
C2664 ALU_1b_2/comparator_0/w_n195_n67# ALU_1b_2/comparator_0/NOR_3/A 0.06fF
C2665 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# ALU_1b_0/full_adder_1/NOR_0/A 0.03fF
C2666 ALU_1b_0/comparator_0/NOR_0/A gnd 0.17fF
C2667 vdd ALU_1b_2/comparator_0/AND_1/w_64_45# 0.14fF
C2668 ALU_1b_2/NOR_0/A ALU_1b_2/AND_5/B 0.01fF
C2669 ALU_1b_2/AND_13/a_78_51# B1 0.19fF
C2670 ALU_1b_2/comparator_0/NOR_2/B ALU_1b_2/AND_11/B 0.10fF
C2671 ALU_1b_0/NOT_5/in ALU_1b_0/NOR_4/B 0.03fF
C2672 ALU_1b_1/AND_17/A ALU_1b_1/full_adder_0/NOR_0/out 0.04fF
C2673 gnd ALU_1b_3/AND_2/a_78_51# 0.07fF
C2674 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.00fF
C2675 ALU_1b_3/AND_18/a_78_51# ALU_1b_3/AND_5/B 0.19fF
C2676 ALU_1b_1/comparator_0/AND_0/w_64_45# ALU_1b_1/comparator_0/AND_2/B 0.06fF
C2677 A2 ALU_1b_3/AND_3/A 0.03fF
C2678 gnd ALU_1b_2/comparator_0/AND_1/a_78_51# 0.07fF
C2679 ALU_1b_3/comparator_0/NOR_2/B ALU_1b_3/comparator_0/NOR_2/out 0.27fF
C2680 ALU_1b_1/AND_14/B B3 0.23fF
C2681 ALU_1b_0/AND_12/a_78_51# vdd 0.06fF
C2682 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/AND_1/out 0.72fF
C2683 ALU_1b_3/AND_10/a_78_51# ALU_1b_3/AND_10/B 0.38fF
C2684 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out ALU_1b_0/full_adder_0/NOR_0/B 0.05fF
C2685 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.05fF
C2686 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# vdd 0.06fF
C2687 ALU_1b_1/AND_5/a_78_51# ALU_1b_1/AND_5/B 0.19fF
C2688 ALU_1b_1/decoder_0/AND_2/B ALU_1b_1/AND_12/w_64_45# 0.06fF
C2689 ALU_1b_0/NOR_2/A vdd 0.03fF
C2690 ALU_1b_0/comparator_0/AND_5/B gnd 0.07fF
C2691 gnd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.14fF
C2692 ALU_1b_1/AND_9/w_64_45# F2 0.06fF
C2693 ALU_1b_2/AND_6/a_78_51# ALU_1b_2/AND_6/out 0.05fF
C2694 S1 ALU_1b_3/decoder_0/AND_2/B 0.07fF
C2695 gnd ALU_1b_3/NOR_0/A 0.17fF
C2696 ALU_1b_2/AND_9/A B1 0.28fF
C2697 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/NOT_1/in 0.23fF
C2698 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/NOR_0/B 0.09fF
C2699 ALU_1b_1/AND_5/w_64_45# vdd 0.15fF
C2700 gnd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.02fF
C2701 ALU_1b_2/AND_0/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.03fF
C2702 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# ALU_1b_3/AND_16/A 0.13fF
C2703 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/A 0.16fF
C2704 vdd ALU_1b_3/AND_5/out 0.35fF
C2705 ALU_1b_0/AND_17/A ALU_1b_0/AND_17/w_64_45# 0.06fF
C2706 ALU_1b_0/decoder_0/AND_1/a_78_51# vdd 0.06fF
C2707 ALU_1b_3/AND_2/out gnd 0.07fF
C2708 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# 0.04fF
C2709 ALU_1b_1/AND_5/a_78_51# gnd 0.07fF
C2710 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# ALU_1b_1/full_adder_1/half_adder_1/A 0.06fF
C2711 ALU_1b_2/comparator_0/w_n220_n67# ALU_1b_2/comparator_0/NOR_2/A 0.06fF
C2712 ALU_1b_0/AND_9/a_78_51# gnd 0.07fF
C2713 A1 ALU_1b_2/AND_12/a_78_51# 0.19fF
C2714 ALU_1b_1/AND_0/a_78_51# ALU_1b_1/AND_0/out 0.05fF
C2715 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C2716 ALU_1b_1/AND_1/a_78_51# ALU_1b_1/AND_2/B 0.19fF
C2717 ALU_1b_1/AND_19/w_64_45# ALU_1b_1/NOR_0/A 0.03fF
C2718 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/comparator_0/AND_5/B 0.17fF
C2719 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/AND_2/a_78_51# 0.19fF
C2720 ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/AND_1/a_78_51# 0.20fF
C2721 S1 ALU_1b_2/C0 0.22fF
C2722 gnd ALU_1b_2/AND_14/A 0.07fF
C2723 ALU_1b_3/AND_9/w_64_45# ALU_1b_3/AND_9/a_78_51# 0.09fF
C2724 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/AND_3/out 0.00fF
C2725 ALU_1b_3/decoder_0/AND_2/B ALU_1b_3/decoder_0/AND_1/B 0.59fF
C2726 ALU_1b_1/decoder_0/AND_2/B gnd 0.07fF
C2727 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/AND_0/out 0.13fF
C2728 ALU_1b_1/NOR_4/w_n27_1# vdd 0.24fF
C2729 vdd ALU_1b_2/comparator_0/NOR_1/B 0.30fF
C2730 ALU_1b_0/AND_8/w_64_45# ALU_1b_0/AND_8/a_78_51# 0.09fF
C2731 ALU_1b_0/AND_11/a_78_51# ALU_1b_0/AND_9/A 0.03fF
C2732 ALU_1b_1/AND_0/out ALU_1b_1/AND_2/B 0.11fF
C2733 vdd ALU_1b_2/AND_15/B 0.09fF
C2734 ALU_1b_0/AND_9/A ALU_1b_0/AND_11/B 0.37fF
C2735 ALU_1b_2/NOT_2/in ALU_1b_2/NOR_2/A 0.03fF
C2736 ALU_1b_3/AND_6/out ALU_1b_3/AND_7/out 0.13fF
C2737 gnd ALU_1b_3/comparator_0/NOR_2/B 0.07fF
C2738 ALU_1b_1/AND_2/out ALU_1b_1/AND_2/a_78_51# 0.05fF
C2739 ALU_1b_1/comparator_0/AND_0/w_64_45# vdd 0.14fF
C2740 ALU_1b_1/comparator_0/AND_3/w_64_45# ALU_1b_1/comparator_0/AND_3/a_78_51# 0.09fF
C2741 ALU_1b_1/AND_9/out ALU_1b_1/AND_7/out 0.02fF
C2742 gnd ALU_1b_2/comparator_0/NOR_1/out 0.07fF
C2743 ALU_1b_1/AND_12/a_78_51# ALU_1b_1/AND_15/A 0.05fF
C2744 vdd ALU_1b_2/AND_1/a_78_51# 0.06fF
C2745 ALU_1b_0/AND_12/w_64_45# ALU_1b_0/decoder_0/AND_1/B 0.03fF
C2746 ALU_1b_1/NOT_3/in gnd 0.07fF
C2747 ALU_1b_2/NOT_1/in ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.13fF
C2748 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_3/B 0.15fF
C2749 ALU_1b_1/comparator_0/AND_0/a_78_51# gnd 0.07fF
C2750 ALU_1b_2/NOR_0/A ALU_1b_2/NOR_3/A 0.01fF
C2751 S1 ALU_1b_1/decoder_0/AND_1/B 0.29fF
C2752 ALU_1b_0/comparator_0/AND_3/w_64_45# ALU_1b_0/AND_8/out 0.16fF
C2753 vdd A2 0.21fF
C2754 ALU_1b_2/AND_9/a_78_51# ALU_1b_2/AND_9/out 0.05fF
C2755 ALU_1b_2/AND_7/a_78_51# ALU_1b_2/AND_8/out 0.10fF
C2756 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/AND_1/out 0.70fF
C2757 ALU_1b_2/comparator_0/w_113_n67# ALU_1b_2/AND_10/B 0.03fF
C2758 ALU_1b_3/AND_18/a_78_51# ALU_1b_3/NOR_3/A 0.07fF
C2759 Cin gnd 0.15fF
C2760 ALU_1b_2/AND_4/w_64_45# B1 0.10fF
C2761 vdd S0 1.80fF
C2762 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out ALU_1b_3/full_adder_1/half_adder_1/A 0.14fF
C2763 ALU_1b_2/AND_0/out vdd 0.03fF
C2764 gnd ALU_1b_2/NOR_3/B 0.23fF
C2765 ALU_1b_1/comparator_0/NOR_0/A ALU_1b_1/comparator_0/NOR_0/out 0.03fF
C2766 ALU_1b_3/NOT_1/in ALU_1b_3/AND_5/out 0.21fF
C2767 ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.10fF
C2768 vdd ALU_1b_2/full_adder_0/NOR_0/out 0.03fF
C2769 vdd ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C2770 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/w_n39_45# 0.11fF
C2771 ALU_1b_0/AND_9/out ALU_1b_0/comparator_0/w_n39_45# 0.15fF
C2772 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out 0.05fF
C2773 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# ALU_1b_0/AND_2/out 0.10fF
C2774 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_0/full_adder_0/NOR_0/B 0.52fF
C2775 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOR_3/A 0.06fF
C2776 ALU_1b_1/AND_15/A vdd 0.43fF
C2777 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.14fF
C2778 ALU_1b_2/AND_4/out ALU_1b_2/AND_5/a_78_51# 0.24fF
C2779 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_15/B 0.03fF
C2780 ALU_1b_1/AND_13/a_78_51# ALU_1b_1/AND_14/B 0.10fF
C2781 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C2782 gnd ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out 0.04fF
C2783 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.06fF
C2784 ALU_1b_2/AND_8/out ALU_1b_2/comparator_0/AND_4/a_78_51# 0.20fF
C2785 ALU_1b_0/AND_3/out ALU_1b_0/AND_5/w_64_45# 0.20fF
C2786 ALU_1b_1/NOR_1/B F2 0.01fF
C2787 ALU_1b_2/AND_15/B ALU_1b_2/AND_15/A 0.28fF
C2788 ALU_1b_0/AND_14/A ALU_1b_0/AND_14/a_78_51# 0.03fF
C2789 ALU_1b_2/AND_6/w_64_45# ALU_1b_2/decoder_0/AND_2/B 0.09fF
C2790 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_10/a_78_51# 0.09fF
C2791 ALU_1b_0/AND_3/a_78_51# ALU_1b_0/AND_5/B 0.29fF
C2792 ALU_1b_1/decoder_0/AND_2/a_78_51# vdd 0.06fF
C2793 ALU_1b_3/AND_1/w_64_45# ALU_1b_3/AND_2/B 0.06fF
C2794 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out 0.20fF
C2795 ALU_1b_3/AND_15/a_78_51# ALU_1b_3/AND_15/A 0.05fF
C2796 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_2/AND_3/out 0.13fF
C2797 ALU_1b_3/AND_18/A ALU_1b_3/AND_5/B 0.26fF
C2798 gnd ALU_1b_2/decoder_0/AND_0/a_78_51# 0.07fF
C2799 vdd ALU_1b_3/comparator_0/w_113_n67# 0.12fF
C2800 ALU_1b_0/comparator_0/w_113_n67# ALU_1b_0/comparator_0/NOR_1/out 0.11fF
C2801 vdd ALU_1b_3/AND_14/a_78_51# 0.06fF
C2802 ALU_1b_1/AND_17/A ALU_1b_1/full_adder_0/w_448_45# 0.03fF
C2803 ALU_1b_0/comparator_0/NOR_3/B gnd 0.21fF
C2804 ALU_1b_3/comparator_0/w_113_n67# ALU_1b_3/comparator_0/NOR_1/B 0.62fF
C2805 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/C0 0.19fF
C2806 vdd ALU_1b_3/AND_0/w_64_45# 0.15fF
C2807 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out 0.05fF
C2808 ALU_1b_3/AND_14/a_78_51# ALU_1b_3/AND_15/B 0.05fF
C2809 ALU_1b_0/AND_5/out C1 0.01fF
C2810 ALU_1b_3/AND_19/A ALU_1b_3/AND_5/B 0.26fF
C2811 gnd ALU_1b_2/AND_6/out 0.07fF
C2812 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_2/a_n14_7# 0.00fF
C2813 vdd ALU_1b_3/AND_17/w_64_45# 0.15fF
C2814 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_74# vdd 0.02fF
C2815 ALU_1b_1/NOR_0/B gnd 0.17fF
C2816 ALU_1b_1/AND_5/out F2 0.01fF
C2817 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/AND_1/out 0.06fF
C2818 vdd ALU_1b_3/comparator_0/w_n74_45# 0.06fF
C2819 ALU_1b_3/AND_16/A ALU_1b_3/AND_16/w_64_45# 0.06fF
C2820 ALU_1b_0/AND_4/out ALU_1b_0/AND_5/a_78_51# 0.24fF
C2821 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_9/out 0.19fF
C2822 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/full_adder_1/half_adder_1/A 0.01fF
C2823 S0 ALU_1b_2/decoder_0/AND_2/a_78_51# 0.05fF
C2824 vdd ALU_1b_2/NOR_2/B 0.03fF
C2825 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/NOR_3/out 0.15fF
C2826 ALU_1b_1/AND_1/out gnd 0.69fF
C2827 gnd ALU_1b_3/AND_17/a_78_51# 0.07fF
C2828 vdd ALU_1b_2/comparator_0/NOR_0/A 0.03fF
C2829 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_0/out 0.23fF
C2830 ALU_1b_2/AND_11/a_78_51# ALU_1b_2/AND_11/B 0.19fF
C2831 ALU_1b_0/AND_4/w_64_45# ALU_1b_0/AND_5/B 0.06fF
C2832 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C2833 ALU_1b_3/AND_8/out B2 0.01fF
C2834 ALU_1b_1/AND_5/B ALU_1b_1/C0 0.28fF
C2835 A3 ALU_1b_1/AND_6/a_78_51# 0.19fF
C2836 vdd B3 0.28fF
C2837 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.00fF
C2838 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/NOR_0/B 0.38fF
C2839 gnd ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C2840 ALU_1b_3/comparator_0/NOR_2/out ALU_1b_3/AND_11/B 0.05fF
C2841 ALU_1b_0/AND_17/w_64_45# ALU_1b_0/NOR_3/B 0.07fF
C2842 ALU_1b_1/AND_6/w_64_45# ALU_1b_1/decoder_0/AND_1/B 0.13fF
C2843 ALU_1b_2/comparator_0/AND_0/w_64_45# ALU_1b_2/comparator_0/NOR_0/A 0.03fF
C2844 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_0/a_78_51# 0.29fF
C2845 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C2846 ALU_1b_3/AND_0/w_64_45# ALU_1b_3/AND_0/out 0.09fF
C2847 ALU_1b_3/full_adder_0/NOR_0/A gnd 0.07fF
C2848 vdd ALU_1b_2/comparator_0/AND_5/B 0.03fF
C2849 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out ALU_1b_3/AND_4/out 0.20fF
C2850 ALU_1b_0/AND_3/A ALU_1b_0/AND_5/B 0.42fF
C2851 ALU_1b_3/AND_6/out ALU_1b_3/AND_9/out 0.29fF
C2852 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/AND_5/B 0.16fF
C2853 gnd ALU_1b_2/comparator_0/NOR_2/A 0.24fF
C2854 ALU_1b_1/AND_9/A ALU_1b_1/AND_6/w_64_45# 0.36fF
C2855 ALU_1b_3/NOR_1/B ALU_1b_3/C0 0.01fF
C2856 ALU_1b_0/AND_7/out vdd 0.34fF
C2857 ALU_1b_1/AND_16/w_64_45# ALU_1b_1/AND_2/B 0.10fF
C2858 ALU_1b_2/AND_19/w_64_45# ALU_1b_2/AND_19/A 0.06fF
C2859 gnd ALU_1b_1/C0 0.69fF
C2860 vdd ALU_1b_3/NOR_4/A 0.10fF
C2861 ALU_1b_1/NOT_1/in ALU_1b_1/AND_18/A 0.12fF
C2862 ALU_1b_2/AND_9/out ALU_1b_2/comparator_0/AND_2/w_64_45# 0.16fF
C2863 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_5/w_64_45# 0.03fF
C2864 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C2865 ALU_1b_0/comparator_0/AND_2/w_64_45# ALU_1b_0/comparator_0/AND_2/a_78_51# 0.09fF
C2866 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_4/w_64_45# 0.03fF
C2867 ALU_1b_0/comparator_0/NOR_3/A ALU_1b_0/AND_7/out 0.11fF
C2868 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/NOR_1/A 0.03fF
C2869 vdd ALU_1b_3/AND_5/a_78_51# 0.06fF
C2870 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.09fF
C2871 vdd ALU_1b_2/AND_9/a_78_51# 0.06fF
C2872 ALU_1b_2/NOR_2/A ALU_1b_2/NOT_3/in 0.23fF
C2873 ALU_1b_1/NOR_0/B ALU_1b_1/NOR_3/A 0.01fF
C2874 ALU_1b_0/full_adder_1/half_adder_1/A gnd 0.03fF
C2875 gnd ALU_1b_2/comparator_0/NOR_0/B 0.17fF
C2876 ALU_1b_2/AND_0/out B1 0.01fF
C2877 ALU_1b_1/NOT_1/in ALU_1b_1/AND_19/A 0.03fF
C2878 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# ALU_1b_1/full_adder_1/half_adder_1/A 0.03fF
C2879 ALU_1b_0/NOR_4/A ALU_1b_0/NOR_1/A 0.01fF
C2880 ALU_1b_2/AND_19/a_78_51# ALU_1b_2/NOR_0/A 0.16fF
C2881 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out 0.09fF
C2882 vdd ALU_1b_3/decoder_0/AND_2/B 0.03fF
C2883 ALU_1b_0/AND_7/a_78_51# ALU_1b_0/AND_7/out 0.16fF
C2884 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_74# vdd 0.02fF
C2885 ALU_1b_0/NOR_1/B gnd 0.22fF
C2886 ALU_1b_0/comparator_0/NOR_3/B ALU_1b_0/comparator_0/AND_4/a_78_8# 0.00fF
C2887 vdd ALU_1b_2/AND_16/w_64_45# 0.15fF
C2888 ALU_1b_3/full_adder_0/half_adder_1/A ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.13fF
C2889 ALU_1b_1/full_adder_1/half_adder_0/w_36_45# ALU_1b_1/AND_4/out 0.29fF
C2890 ALU_1b_2/AND_5/w_64_45# ALU_1b_2/C0 0.10fF
C2891 gnd ALU_1b_3/AND_11/a_78_51# 0.07fF
C2892 vdd ALU_1b_2/full_adder_0/w_448_45# 0.12fF
C2893 ALU_1b_3/AND_7/w_64_45# ALU_1b_3/AND_7/out 0.03fF
C2894 ALU_1b_3/AND_5/out ALU_1b_3/C0 0.01fF
C2895 gnd ALU_1b_3/AND_11/B 0.13fF
C2896 gnd ALU_1b_2/AND_16/a_78_51# 0.07fF
C2897 ALU_1b_2/AND_12/w_64_45# ALU_1b_2/AND_5/B 0.03fF
C2898 ALU_1b_0/AND_16/A ALU_1b_0/AND_2/B 0.26fF
C2899 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C2900 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.09fF
C2901 ALU_1b_1/AND_9/A ALU_1b_1/AND_10/B 0.29fF
C2902 ALU_1b_1/NOR_4/A ALU_1b_1/AND_11/a_78_51# 0.07fF
C2903 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C2904 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C2905 vdd ALU_1b_3/comparator_0/AND_0/a_78_51# 0.06fF
C2906 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/w_n74_45# 0.18fF
C2907 ALU_1b_0/AND_12/a_78_51# ALU_1b_0/AND_14/B 0.05fF
C2908 ALU_1b_1/AND_1/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.05fF
C2909 ALU_1b_2/AND_3/a_78_51# ALU_1b_2/AND_3/A 0.03fF
C2910 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.06fF
C2911 ALU_1b_0/AND_5/out vdd 0.35fF
C2912 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# gnd 0.14fF
C2913 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_74# 0.01fF
C2914 ALU_1b_3/AND_4/out ALU_1b_3/full_adder_1/half_adder_1/A 0.11fF
C2915 ALU_1b_2/NOR_2/A ALU_1b_2/NOR_2/w_n27_1# 0.06fF
C2916 vdd ALU_1b_2/C0 0.56fF
C2917 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.00fF
C2918 ALU_1b_1/comparator_0/AND_3/a_78_51# ALU_1b_1/AND_8/out 0.03fF
C2919 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/comparator_0/AND_4/a_78_51# 0.04fF
C2920 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_1/half_adder_1/A 0.13fF
C2921 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out vdd 0.06fF
C2922 ALU_1b_0/full_adder_1/NOR_0/A gnd 0.07fF
C2923 ALU_1b_3/AND_14/B ALU_1b_3/AND_12/w_64_45# 0.03fF
C2924 gnd ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.04fF
C2925 vdd ALU_1b_3/comparator_0/AND_3/w_64_45# 0.15fF
C2926 ALU_1b_1/comparator_0/NOR_1/A gnd 0.17fF
C2927 ALU_1b_3/AND_4/a_78_51# B2 0.03fF
C2928 ALU_1b_1/decoder_0/AND_1/a_78_51# ALU_1b_1/decoder_0/AND_1/B 0.19fF
C2929 ALU_1b_0/AND_7/out ALU_1b_0/comparator_0/AND_4/a_78_51# 0.03fF
C2930 ALU_1b_2/AND_14/w_64_45# ALU_1b_2/AND_14/A 0.09fF
C2931 ALU_1b_1/AND_4/out ALU_1b_1/AND_4/w_64_45# 0.03fF
C2932 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_1/AND_3/out 0.03fF
C2933 ALU_1b_3/NOR_4/w_n27_1# ALU_1b_3/NOR_3/B 0.20fF
C2934 ALU_1b_0/AND_3/out B0 0.01fF
C2935 vdd ALU_1b_3/AND_2/w_64_45# 0.15fF
C2936 ALU_1b_3/comparator_0/AND_4/w_64_45# ALU_1b_3/AND_7/out 0.10fF
C2937 gnd ALU_1b_3/comparator_0/AND_3/a_78_51# 0.07fF
C2938 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C2939 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_0/half_adder_1/A 0.26fF
C2940 ALU_1b_3/AND_14/A ALU_1b_3/AND_15/A 0.10fF
C2941 ALU_1b_2/decoder_0/AND_0/a_78_51# ALU_1b_2/AND_2/B 0.05fF
C2942 ALU_1b_1/NOT_5/in ALU_1b_1/NOR_4/w_n27_1# 0.11fF
C2943 ALU_1b_1/AND_13/a_78_51# vdd 0.06fF
C2944 gnd ALU_1b_3/AND_5/B 0.48fF
C2945 ALU_1b_1/decoder_0/AND_1/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C2946 ALU_1b_1/AND_3/out ALU_1b_1/AND_5/out 0.11fF
C2947 ALU_1b_0/AND_2/out C1 0.01fF
C2948 ALU_1b_1/AND_8/out gnd 0.23fF
C2949 vdd ALU_1b_1/decoder_0/AND_1/B 0.03fF
C2950 ALU_1b_0/comparator_0/NOR_0/B ALU_1b_0/comparator_0/w_113_n67# 0.02fF
C2951 ALU_1b_0/comparator_0/w_88_n67# ALU_1b_0/comparator_0/NOR_1/B 0.19fF
C2952 ALU_1b_1/full_adder_1/NOR_0/B gnd 0.07fF
C2953 vdd ALU_1b_3/NOR_2/w_n27_1# 0.24fF
C2954 ALU_1b_0/AND_0/w_64_45# ALU_1b_0/AND_2/B 0.06fF
C2955 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out ALU_1b_2/full_adder_1/NOR_0/B 0.00fF
C2956 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_1/AND_1/out 0.10fF
C2957 vdd ALU_1b_2/AND_9/w_64_45# 0.42fF
C2958 C0 Cin 3.17fF
C2959 ALU_1b_3/AND_8/out ALU_1b_3/AND_9/A 0.12fF
C2960 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/w_n74_45# 0.03fF
C2961 ALU_1b_0/decoder_0/AND_0/a_78_51# ALU_1b_0/decoder_0/AND_2/B 0.03fF
C2962 ALU_1b_1/AND_15/w_64_45# vdd 0.15fF
C2963 ALU_1b_1/AND_9/A vdd 1.07fF
C2964 ALU_1b_1/AND_19/w_64_45# ALU_1b_1/AND_5/B 0.06fF
C2965 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/NOT_1/in 0.06fF
C2966 gnd ALU_1b_2/AND_10/a_78_51# 0.07fF
C2967 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.06fF
C2968 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_0/NOT_1/in 0.06fF
C2969 ALU_1b_1/AND_15/a_78_51# gnd 0.07fF
C2970 ALU_1b_2/comparator_0/NOR_0/B ALU_1b_2/comparator_0/NOR_0/out 0.15fF
C2971 ALU_1b_2/AND_7/out ALU_1b_2/comparator_0/w_n74_45# 0.10fF
C2972 ALU_1b_3/AND_0/out ALU_1b_3/AND_2/w_64_45# 0.20fF
C2973 ALU_1b_1/NOR_4/A gnd 0.23fF
C2974 ALU_1b_2/AND_15/B ALU_1b_2/AND_15/w_64_45# 0.06fF
C2975 ALU_1b_2/NOR_1/B ALU_1b_2/NOR_1/A 0.33fF
C2976 ALU_1b_2/comparator_0/w_n220_n67# ALU_1b_2/comparator_0/NOR_2/B 0.62fF
C2977 A0 gnd 0.48fF
C2978 ALU_1b_2/full_adder_0/NOR_0/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.06fF
C2979 vdd ALU_1b_2/comparator_0/NOR_3/B 0.03fF
C2980 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/AND_0/out 0.10fF
C2981 ALU_1b_1/AND_1/w_64_45# vdd 0.15fF
C2982 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/a_n7_n34# ALU_1b_1/AND_1/out 0.00fF
C2983 ALU_1b_3/AND_15/w_64_45# ALU_1b_3/AND_15/a_78_51# 0.09fF
C2984 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/NOR_0/out 0.15fF
C2985 ALU_1b_0/AND_0/w_64_45# vdd 0.15fF
C2986 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# ALU_1b_3/AND_5/out 0.10fF
C2987 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# vdd 0.22fF
C2988 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.00fF
C2989 ALU_1b_1/AND_3/a_78_51# vdd 0.06fF
C2990 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_2/full_adder_1/half_adder_1/A 0.13fF
C2991 S0 ALU_1b_2/decoder_0/AND_1/B 0.03fF
C2992 ALU_1b_1/comparator_0/NOR_3/A ALU_1b_1/comparator_0/NOR_3/B 0.43fF
C2993 gnd ALU_1b_2/comparator_0/NOR_3/out 0.07fF
C2994 ALU_1b_0/AND_9/out vdd 0.86fF
C2995 ALU_1b_0/decoder_0/AND_2/a_78_51# S1 0.02fF
C2996 ALU_1b_1/AND_7/out B3 0.28fF
C2997 ALU_1b_0/AND_0/a_78_51# gnd 0.07fF
C2998 ALU_1b_1/full_adder_1/half_adder_0/w_36_45# vdd 0.14fF
C2999 vdd ALU_1b_3/NOR_0/B 0.20fF
C3000 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out ALU_1b_0/AND_5/out 0.08fF
C3001 ALU_1b_2/full_adder_1/NOR_0/A ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C3002 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_0/a_78_51# 0.14fF
C3003 ALU_1b_0/decoder_0/AND_1/a_78_51# ALU_1b_0/AND_6/w_64_45# 0.09fF
C3004 ALU_1b_0/NOT_2/in gnd 0.07fF
C3005 vdd ALU_1b_2/comparator_0/AND_2/w_64_45# 0.15fF
C3006 vdd ALU_1b_3/AND_1/out 0.35fF
C3007 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C3008 ALU_1b_3/comparator_0/AND_0/w_64_45# ALU_1b_3/AND_6/out 0.26fF
C3009 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_36# ALU_1b_3/AND_16/A 0.03fF
C3010 ALU_1b_1/comparator_0/AND_0/w_64_45# ALU_1b_1/AND_9/out 0.30fF
C3011 gnd ALU_1b_2/comparator_0/AND_2/a_78_51# 0.07fF
C3012 ALU_1b_0/AND_0/out gnd 0.11fF
C3013 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.09fF
C3014 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# gnd 0.02fF
C3015 ALU_1b_1/full_adder_0/NOR_0/A ALU_1b_1/AND_1/out 0.04fF
C3016 ALU_1b_0/AND_8/a_78_51# vdd 0.06fF
C3017 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/AND_5/out 0.02fF
C3018 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# ALU_1b_2/AND_1/out 0.29fF
C3019 ALU_1b_1/AND_4/a_78_51# ALU_1b_1/AND_5/B 0.29fF
C3020 ALU_1b_0/AND_2/out ALU_1b_0/AND_2/B 0.38fF
C3021 ALU_1b_2/AND_8/out ALU_1b_2/AND_6/w_64_45# 0.15fF
C3022 ALU_1b_3/AND_4/out ALU_1b_3/AND_5/B 0.38fF
C3023 gnd ALU_1b_3/NOR_3/A 0.23fF
C3024 vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.06fF
C3025 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_74# vdd 0.02fF
C3026 ALU_1b_3/AND_1/out ALU_1b_3/AND_1/a_78_51# 0.05fF
C3027 ALU_1b_3/NOT_3/in ALU_1b_3/NOR_2/B 0.03fF
C3028 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_0/full_adder_0/half_adder_1/A 0.13fF
C3029 ALU_1b_1/AND_17/a_78_51# ALU_1b_1/NOR_3/B 0.07fF
C3030 ALU_1b_1/AND_16/A ALU_1b_1/AND_2/B 0.26fF
C3031 ALU_1b_3/comparator_0/AND_0/a_78_51# ALU_1b_3/comparator_0/NOR_0/A 0.05fF
C3032 ALU_1b_3/NOT_6/in ALU_1b_3/NOR_4/B 0.15fF
C3033 ALU_1b_1/AND_4/w_64_45# vdd 0.15fF
C3034 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_2/A 0.33fF
C3035 ALU_1b_1/AND_2/out gnd 0.07fF
C3036 ALU_1b_2/full_adder_1/NOR_0/A vdd 0.03fF
C3037 ALU_1b_0/NOR_1/A vdd 0.22fF
C3038 ALU_1b_3/full_adder_0/NOR_0/A ALU_1b_3/full_adder_0/half_adder_1/w_36_45# 0.03fF
C3039 ALU_1b_1/AND_4/a_78_51# gnd 0.07fF
C3040 ALU_1b_2/NOT_4/in ALU_1b_2/NOR_2/w_n27_1# 0.11fF
C3041 ALU_1b_0/AND_14/a_78_51# gnd 0.07fF
C3042 ALU_1b_3/AND_1/out ALU_1b_3/AND_0/out 0.11fF
C3043 ALU_1b_0/decoder_0/AND_3/a_78_51# ALU_1b_0/AND_15/A 0.05fF
C3044 ALU_1b_3/full_adder_0/NOR_0/B ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.00fF
C3045 ALU_1b_1/NOR_4/w_n27_1# ALU_1b_1/NOR_1/A 0.09fF
C3046 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_3/full_adder_1/half_adder_1/A 0.03fF
C3047 ALU_1b_1/AND_3/w_64_45# A3 0.10fF
C3048 ALU_1b_2/AND_16/a_78_51# ALU_1b_2/AND_2/B 0.19fF
C3049 ALU_1b_3/AND_3/out ALU_1b_3/AND_3/w_64_45# 0.09fF
C3050 ALU_1b_3/AND_19/A ALU_1b_3/AND_19/a_78_51# 0.03fF
C3051 ALU_1b_0/AND_2/out vdd 0.35fF
C3052 ALU_1b_0/full_adder_1/NOR_0/out ALU_1b_0/NOT_1/in 0.10fF
C3053 ALU_1b_3/AND_1/out ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# 0.06fF
C3054 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_16/A 0.23fF
C3055 ALU_1b_3/comparator_0/NOR_3/A ALU_1b_3/comparator_0/AND_5/a_78_51# 0.05fF
C3056 ALU_1b_3/AND_9/out ALU_1b_3/comparator_0/AND_2/a_78_51# 0.03fF
C3057 ALU_1b_2/C0 B1 2.34fF
C3058 gnd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.11fF
C3059 ALU_1b_1/comparator_0/NOR_3/B ALU_1b_1/comparator_0/AND_4/a_78_51# 0.18fF
C3060 ALU_1b_1/AND_3/A vdd 0.03fF
C3061 ALU_1b_1/NOT_2/in ALU_1b_1/NOR_0/w_n27_1# 0.11fF
C3062 ALU_1b_3/AND_10/a_78_51# ALU_1b_3/NOR_1/A 0.05fF
C3063 ALU_1b_3/AND_3/out F1 0.01fF
C3064 ALU_1b_0/full_adder_0/NOR_0/B gnd 0.07fF
C3065 ALU_1b_2/AND_18/w_64_45# ALU_1b_2/AND_18/a_78_51# 0.09fF
C3066 ALU_1b_3/AND_12/a_78_51# ALU_1b_3/AND_12/w_64_45# 0.09fF
C3067 vdd ALU_1b_3/comparator_0/w_n195_n67# 0.12fF
C3068 ALU_1b_0/comparator_0/AND_3/w_64_45# ALU_1b_0/comparator_0/NOR_2/A 0.03fF
C3069 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_3/a_78_51# 0.19fF
C3070 ALU_1b_0/comparator_0/NOR_0/A ALU_1b_0/comparator_0/w_88_n67# 0.06fF
C3071 ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# 0.26fF
C3072 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_74# ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.01fF
C3073 ALU_1b_0/AND_6/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C3074 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# 0.13fF
C3075 vdd ALU_1b_2/NOR_1/B 0.20fF
C3076 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/A 0.06fF
C3077 ALU_1b_2/AND_5/out ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.06fF
C3078 ALU_1b_3/comparator_0/AND_3/w_64_45# ALU_1b_3/comparator_0/AND_5/B 0.06fF
C3079 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_0/AND_1/out 0.10fF
C3080 ALU_1b_1/comparator_0/AND_1/w_64_45# vdd 0.14fF
C3081 ALU_1b_3/NOR_2/B ALU_1b_3/NOR_2/w_n27_1# 0.09fF
C3082 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# ALU_1b_3/AND_5/out 0.04fF
C3083 gnd ALU_1b_2/AND_2/a_78_51# 0.07fF
C3084 ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/AND_10/B 0.09fF
C3085 ALU_1b_0/AND_3/out ALU_1b_0/AND_3/a_78_51# 0.05fF
C3086 ALU_1b_1/comparator_0/AND_1/a_78_51# gnd 0.07fF
C3087 ALU_1b_3/AND_5/a_78_51# ALU_1b_3/C0 0.03fF
C3088 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out vdd 0.06fF
C3089 ALU_1b_0/comparator_0/AND_5/w_64_45# ALU_1b_0/AND_8/out 0.32fF
C3090 ALU_1b_2/AND_5/out ALU_1b_2/AND_5/w_64_45# 0.03fF
C3091 ALU_1b_0/AND_8/w_64_45# ALU_1b_0/AND_9/A 0.39fF
C3092 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# 0.03fF
C3093 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# ALU_1b_3/full_adder_0/NOR_0/B 0.00fF
C3094 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# gnd 0.14fF
C3095 S1 ALU_1b_2/decoder_0/AND_2/B 0.07fF
C3096 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/full_adder_1/half_adder_0/w_36_45# 0.12fF
C3097 gnd ALU_1b_2/NOR_0/A 0.17fF
C3098 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/w_36_45# 0.29fF
C3099 ALU_1b_0/AND_16/A ALU_1b_0/full_adder_0/NOR_0/A 0.22fF
C3100 gnd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# 0.14fF
C3101 ALU_1b_3/AND_2/out ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out 0.20fF
C3102 ALU_1b_0/AND_5/w_64_45# vdd 0.15fF
C3103 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# gnd 0.02fF
C3104 vdd ALU_1b_3/comparator_0/NOR_1/A 0.03fF
C3105 ALU_1b_0/AND_0/out ALU_1b_0/AND_2/w_64_45# 0.20fF
C3106 ALU_1b_1/AND_0/a_78_51# A3 0.19fF
C3107 ALU_1b_2/AND_3/out ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.26fF
C3108 ALU_1b_0/comparator_0/NOR_1/A ALU_1b_0/comparator_0/NOR_1/out 0.03fF
C3109 vdd ALU_1b_2/AND_5/out 0.35fF
C3110 C0 ALU_1b_0/NOR_1/B 0.01fF
C3111 ALU_1b_2/AND_2/out gnd 0.07fF
C3112 ALU_1b_0/AND_5/a_78_51# gnd 0.07fF
C3113 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# ALU_1b_0/full_adder_1/NOR_0/B 0.00fF
C3114 ALU_1b_3/comparator_0/NOR_1/A ALU_1b_3/comparator_0/NOR_1/B 0.33fF
C3115 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C3116 ALU_1b_3/NOR_4/A ALU_1b_3/AND_9/w_64_45# 0.03fF
C3117 ALU_1b_1/AND_7/out ALU_1b_1/AND_9/A 0.01fF
C3118 ALU_1b_3/AND_13/a_78_51# ALU_1b_3/AND_14/A 0.05fF
C3119 ALU_1b_2/AND_4/out ALU_1b_2/AND_4/a_78_51# 0.05fF
C3120 ALU_1b_3/full_adder_0/half_adder_1/w_36_45# ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out 0.09fF
C3121 ALU_1b_1/AND_2/out ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# 0.06fF
C3122 ALU_1b_0/AND_0/out ALU_1b_0/AND_2/a_78_51# 0.10fF
C3123 ALU_1b_3/AND_4/w_64_45# ALU_1b_3/AND_4/a_78_51# 0.09fF
C3124 ALU_1b_2/full_adder_0/NOR_0/B ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.52fF
C3125 ALU_1b_1/AND_14/A gnd 0.07fF
C3126 vdd ALU_1b_3/AND_8/out 0.66fF
C3127 ALU_1b_1/AND_3/out ALU_1b_1/AND_5/a_78_51# 0.10fF
C3128 ALU_1b_0/AND_3/out ALU_1b_0/AND_4/w_64_45# 0.20fF
C3129 A3 ALU_1b_1/AND_2/B 0.50fF
C3130 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/AND_4/out 0.09fF
C3131 ALU_1b_2/AND_14/A ALU_1b_2/AND_14/B 0.42fF
C3132 ALU_1b_2/AND_9/a_78_51# ALU_1b_2/AND_9/A 0.05fF
C3133 ALU_1b_0/NOR_0/A ALU_1b_0/NOT_2/in 0.03fF
C3134 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/full_adder_0/w_448_45# 0.16fF
C3135 ALU_1b_0/decoder_0/AND_2/B gnd 0.07fF
C3136 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_11/a_78_51# 0.09fF
C3137 ALU_1b_1/NOT_1/in ALU_1b_1/full_adder_1/NOR_0/out 0.10fF
C3138 ALU_1b_0/AND_9/w_64_45# ALU_1b_0/AND_11/B 0.11fF
C3139 vdd ALU_1b_1/comparator_0/NOR_1/B 0.30fF
C3140 ALU_1b_1/AND_1/out F2 0.01fF
C3141 ALU_1b_1/AND_15/B vdd 0.09fF
C3142 Cin ALU_1b_0/AND_5/B 0.27fF
C3143 ALU_1b_1/full_adder_0/half_adder_1/A ALU_1b_1/AND_16/A 0.23fF
C3144 gnd ALU_1b_2/comparator_0/NOR_2/B 0.07fF
C3145 ALU_1b_0/comparator_0/AND_0/w_64_45# vdd 0.14fF
C3146 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.03fF
C3147 ALU_1b_1/comparator_0/NOR_1/out gnd 0.07fF
C3148 ALU_1b_1/AND_17/A ALU_1b_1/AND_17/w_64_45# 0.06fF
C3149 ALU_1b_2/NOR_0/A ALU_1b_2/NOR_0/w_n27_1# 0.06fF
C3150 vdd ALU_1b_3/AND_15/a_78_51# 0.06fF
C3151 ALU_1b_1/AND_1/a_78_51# vdd 0.06fF
C3152 ALU_1b_0/NOT_3/in gnd 0.07fF
C3153 ALU_1b_0/comparator_0/AND_0/a_78_51# gnd 0.07fF
C3154 ALU_1b_2/AND_19/a_78_51# ALU_1b_2/AND_5/B 0.19fF
C3155 ALU_1b_0/decoder_0/AND_1/B S1 0.29fF
C3156 ALU_1b_2/comparator_0/w_n220_n67# ALU_1b_2/AND_11/B 0.03fF
C3157 ALU_1b_0/NOR_4/w_n27_1# ALU_1b_0/NOR_4/A 0.10fF
C3158 vdd A1 0.21fF
C3159 ALU_1b_3/AND_15/B ALU_1b_3/AND_15/a_78_51# 0.19fF
C3160 vdd ALU_1b_3/full_adder_1/half_adder_1/w_36_45# 0.14fF
C3161 ALU_1b_0/full_adder_1/w_448_45# ALU_1b_0/full_adder_1/NOR_0/B 0.16fF
C3162 ALU_1b_1/AND_8/w_64_45# ALU_1b_1/C0 0.06fF
C3163 ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# 0.26fF
C3164 ALU_1b_3/comparator_0/w_n220_n67# ALU_1b_3/comparator_0/NOR_2/out 0.11fF
C3165 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/comparator_0/NOR_3/out 0.05fF
C3166 gnd ALU_1b_3/NOT_6/in 0.07fF
C3167 ALU_1b_1/AND_0/out vdd 0.03fF
C3168 vdd ALU_1b_3/AND_19/w_64_45# 0.15fF
C3169 ALU_1b_1/NOR_3/B gnd 0.23fF
C3170 ALU_1b_0/full_adder_0/half_adder_1/A ALU_1b_0/AND_2/out 0.11fF
C3171 ALU_1b_0/AND_1/out ALU_1b_0/AND_0/out 0.11fF
C3172 ALU_1b_1/full_adder_0/NOR_0/out vdd 0.03fF
C3173 ALU_1b_0/AND_16/a_78_51# ALU_1b_0/NOR_0/B 0.05fF
C3174 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# vdd 0.06fF
C3175 ALU_1b_1/C0 F2 11.26fF
C3176 ALU_1b_1/NOR_4/A ALU_1b_1/NOT_6/in 0.03fF
C3177 ALU_1b_0/AND_4/out ALU_1b_0/AND_4/a_78_51# 0.05fF
C3178 ALU_1b_0/AND_7/out ALU_1b_0/AND_6/w_64_45# 0.13fF
C3179 ALU_1b_2/full_adder_1/NOR_0/B ALU_1b_2/full_adder_1/NOR_0/out 0.15fF
C3180 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/NOR_3/out 0.03fF
C3181 S1 ALU_1b_3/decoder_0/AND_0/a_78_51# 0.02fF
C3182 gnd ALU_1b_3/AND_19/a_78_51# 0.07fF
C3183 ALU_1b_2/AND_9/A ALU_1b_2/C0 0.28fF
C3184 ALU_1b_1/AND_0/w_64_45# ALU_1b_1/AND_0/a_78_51# 0.09fF
C3185 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_1/AND_16/A 0.06fF
C3186 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.01fF
C3187 ALU_1b_3/AND_16/w_64_45# ALU_1b_3/NOR_0/B 0.03fF
C3188 ALU_1b_0/NOR_2/A ALU_1b_0/NOT_4/in 0.03fF
C3189 ALU_1b_2/full_adder_1/w_448_45# ALU_1b_2/AND_18/A 0.03fF
C3190 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_1/half_adder_1/A 0.03fF
C3191 ALU_1b_2/AND_2/out F0 0.01fF
C3192 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/NOR_0/A 0.12fF
C3193 ALU_1b_0/AND_3/out ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# 0.03fF
C3194 ALU_1b_0/AND_15/A vdd 0.43fF
C3195 F1 ALU_1b_3/AND_2/B 0.01fF
C3196 ALU_1b_2/AND_0/out ALU_1b_2/AND_1/a_78_51# 0.10fF
C3197 ALU_1b_2/AND_18/A ALU_1b_2/AND_18/w_64_45# 0.06fF
C3198 ALU_1b_2/NOR_4/A ALU_1b_2/NOR_1/A 0.01fF
C3199 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# ALU_1b_3/AND_4/out 0.06fF
C3200 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out gnd 0.04fF
C3201 ALU_1b_2/comparator_0/AND_0/a_78_51# ALU_1b_2/AND_9/out 0.02fF
C3202 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/AND_1/a_78_51# 0.10fF
C3203 ALU_1b_3/AND_17/A ALU_1b_3/AND_2/B 0.26fF
C3204 ALU_1b_2/AND_7/w_64_45# ALU_1b_2/AND_7/a_78_51# 0.09fF
C3205 ALU_1b_1/AND_0/w_64_45# ALU_1b_1/AND_2/B 0.06fF
C3206 ALU_1b_2/NOR_1/B B1 0.01fF
C3207 ALU_1b_1/AND_19/w_64_45# ALU_1b_1/AND_19/a_78_51# 0.09fF
C3208 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/full_adder_0/half_adder_1/A 0.14fF
C3209 ALU_1b_3/comparator_0/AND_1/w_64_45# ALU_1b_3/comparator_0/AND_1/a_78_51# 0.09fF
C3210 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.09fF
C3211 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out ALU_1b_2/AND_3/out 0.14fF
C3212 ALU_1b_0/decoder_0/AND_2/a_78_51# vdd 0.06fF
C3213 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# ALU_1b_0/full_adder_1/NOR_0/B 0.00fF
C3214 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.01fF
C3215 ALU_1b_1/AND_17/w_64_45# ALU_1b_1/AND_2/B 0.06fF
C3216 ALU_1b_1/NOR_2/A ALU_1b_1/NOR_2/B 0.47fF
C3217 ALU_1b_3/decoder_0/AND_0/a_78_51# ALU_1b_3/decoder_0/AND_1/B 0.29fF
C3218 ALU_1b_0/AND_1/out ALU_1b_0/full_adder_0/NOR_0/B 0.06fF
C3219 ALU_1b_1/decoder_0/AND_0/a_78_51# gnd 0.07fF
C3220 ALU_1b_3/AND_1/out ALU_1b_3/C0 0.01fF
C3221 ALU_1b_0/AND_6/out ALU_1b_0/AND_8/out 0.10fF
C3222 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/AND_7/out 0.05fF
C3223 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.09fF
C3224 ALU_1b_2/AND_9/w_64_45# ALU_1b_2/AND_9/A 0.95fF
C3225 A1 ALU_1b_2/AND_15/A 0.42fF
C3226 vdd ALU_1b_2/comparator_0/w_113_n67# 0.12fF
C3227 vdd ALU_1b_3/AND_4/a_78_51# 0.06fF
C3228 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# ALU_1b_1/NOT_1/in 0.03fF
C3229 ALU_1b_2/comparator_0/NOR_2/out ALU_1b_2/comparator_0/NOR_2/A 0.03fF
C3230 vdd ALU_1b_2/AND_14/a_78_51# 0.06fF
C3231 ALU_1b_2/AND_2/a_78_51# ALU_1b_2/AND_2/B 0.29fF
C3232 ALU_1b_1/NOR_3/B ALU_1b_1/NOR_3/A 0.34fF
C3233 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# ALU_1b_0/AND_1/out 0.29fF
C3234 ALU_1b_1/AND_6/a_78_51# ALU_1b_1/AND_8/out 0.11fF
C3235 ALU_1b_2/AND_0/w_64_45# vdd 0.15fF
C3236 vdd ALU_1b_3/full_adder_1/NOR_0/B 0.91fF
C3237 B0 ALU_1b_0/AND_2/B 0.28fF
C3238 ALU_1b_0/AND_0/out C0 0.01fF
C3239 ALU_1b_1/AND_6/out gnd 0.07fF
C3240 ALU_1b_2/NOR_1/A ALU_1b_2/NOT_3/in 0.03fF
C3241 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_74# 0.01fF
C3242 ALU_1b_2/comparator_0/NOR_3/A ALU_1b_2/comparator_0/AND_4/a_78_8# 0.00fF
C3243 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_15/A 0.50fF
C3244 ALU_1b_0/NOR_0/B gnd 0.17fF
C3245 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_36# ALU_1b_2/NOT_1/in 0.03fF
C3246 vdd ALU_1b_2/AND_17/w_64_45# 0.15fF
C3247 ALU_1b_3/AND_0/a_78_51# ALU_1b_3/AND_2/B 0.14fF
C3248 vdd ALU_1b_2/comparator_0/w_n74_45# 0.06fF
C3249 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out 0.08fF
C3250 gnd ALU_1b_3/AND_6/a_78_51# 0.07fF
C3251 ALU_1b_1/decoder_0/AND_2/a_78_51# S0 0.05fF
C3252 vdd ALU_1b_1/NOR_2/B 0.03fF
C3253 ALU_1b_3/AND_6/out ALU_1b_3/AND_9/A 0.01fF
C3254 ALU_1b_1/AND_8/w_64_45# ALU_1b_1/AND_8/out 0.03fF
C3255 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out ALU_1b_0/full_adder_0/NOR_0/A 0.05fF
C3256 ALU_1b_1/comparator_0/NOR_0/A vdd 0.03fF
C3257 ALU_1b_1/comparator_0/AND_3/a_78_51# ALU_1b_1/comparator_0/NOR_2/A 0.17fF
C3258 ALU_1b_1/AND_9/out ALU_1b_1/AND_9/A 0.04fF
C3259 gnd ALU_1b_2/AND_17/a_78_51# 0.07fF
C3260 ALU_1b_2/AND_2/out ALU_1b_2/AND_2/B 0.38fF
C3261 ALU_1b_3/AND_0/w_64_45# A2 0.10fF
C3262 vdd ALU_1b_3/comparator_0/AND_1/a_78_51# 0.06fF
C3263 B0 vdd 0.28fF
C3264 ALU_1b_2/full_adder_1/half_adder_1/A gnd 0.03fF
C3265 ALU_1b_2/comparator_0/NOR_1/out ALU_1b_2/AND_10/B 0.05fF
C3266 ALU_1b_2/AND_5/w_64_45# ALU_1b_2/AND_5/a_78_51# 0.09fF
C3267 ALU_1b_3/NOR_1/B ALU_1b_3/NOT_3/in 0.15fF
C3268 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/AND_8/out 0.38fF
C3269 ALU_1b_2/full_adder_0/NOR_0/A gnd 0.07fF
C3270 ALU_1b_1/comparator_0/AND_5/a_78_51# ALU_1b_1/AND_8/out 0.02fF
C3271 ALU_1b_1/comparator_0/AND_5/B vdd 0.03fF
C3272 ALU_1b_3/AND_5/out ALU_1b_3/AND_5/a_78_51# 0.05fF
C3273 ALU_1b_1/AND_14/w_64_45# ALU_1b_1/AND_14/a_78_51# 0.09fF
C3274 ALU_1b_1/AND_8/a_78_51# ALU_1b_1/AND_9/A 0.05fF
C3275 ALU_1b_0/NOR_2/w_n27_1# F0 0.03fF
C3276 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# ALU_1b_2/AND_4/out 0.70fF
C3277 ALU_1b_2/AND_3/out ALU_1b_2/full_adder_1/half_adder_1/A 0.23fF
C3278 vdd ALU_1b_3/comparator_0/AND_5/w_64_45# 0.13fF
C3279 ALU_1b_1/comparator_0/NOR_2/A gnd 0.24fF
C3280 ALU_1b_2/comparator_0/AND_4/w_64_45# ALU_1b_2/comparator_0/AND_4/a_78_51# 0.09fF
C3281 ALU_1b_2/AND_7/out ALU_1b_2/AND_8/out 0.40fF
C3282 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_74# ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.01fF
C3283 ALU_1b_2/AND_14/a_78_51# ALU_1b_2/AND_15/A 0.00fF
C3284 C1 ALU_1b_0/AND_9/A 0.28fF
C3285 ALU_1b_2/NOR_4/A vdd 0.10fF
C3286 ALU_1b_2/NOR_1/A ALU_1b_2/NOR_2/w_n27_1# 0.10fF
C3287 ALU_1b_2/AND_6/w_64_45# ALU_1b_2/decoder_0/AND_0/a_78_51# 0.09fF
C3288 gnd ALU_1b_3/comparator_0/AND_5/a_78_51# 0.07fF
C3289 ALU_1b_1/comparator_0/w_88_n67# ALU_1b_1/comparator_0/NOR_0/B 0.20fF
C3290 A1 B1 0.65fF
C3291 vdd ALU_1b_2/AND_5/a_78_51# 0.06fF
C3292 ALU_1b_3/full_adder_1/NOR_0/B ALU_1b_3/NOT_1/in 0.06fF
C3293 ALU_1b_0/AND_7/a_78_51# B0 0.19fF
C3294 ALU_1b_1/AND_9/a_78_51# vdd 0.06fF
C3295 ALU_1b_1/NOR_0/B ALU_1b_1/NOR_0/w_n27_1# 0.06fF
C3296 ALU_1b_2/NOR_4/A ALU_1b_2/NOR_4/w_n27_1# 0.10fF
C3297 ALU_1b_1/NOR_1/A ALU_1b_1/AND_9/A 0.03fF
C3298 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_74# ALU_1b_1/AND_16/A 0.03fF
C3299 ALU_1b_1/full_adder_0/NOR_0/B ALU_1b_1/AND_16/A 0.05fF
C3300 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/a_n7_n34# ALU_1b_3/AND_5/out 0.00fF
C3301 ALU_1b_1/AND_3/out ALU_1b_1/C0 0.01fF
C3302 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# ALU_1b_0/AND_0/out 0.09fF
C3303 ALU_1b_1/comparator_0/NOR_0/B gnd 0.17fF
C3304 ALU_1b_3/AND_7/w_64_45# B2 0.06fF
C3305 vdd ALU_1b_3/AND_14/A 0.03fF
C3306 ALU_1b_2/AND_6/out ALU_1b_2/AND_6/w_64_45# 0.14fF
C3307 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_3/AND_5/out 0.70fF
C3308 ALU_1b_0/NOR_4/w_n27_1# vdd 0.24fF
C3309 vdd ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.22fF
C3310 ALU_1b_0/AND_14/w_64_45# B0 0.06fF
C3311 ALU_1b_1/AND_16/w_64_45# vdd 0.15fF
C3312 vdd ALU_1b_2/decoder_0/AND_2/B 0.03fF
C3313 ALU_1b_3/NOR_1/B ALU_1b_3/NOR_2/w_n27_1# 0.06fF
C3314 ALU_1b_1/AND_18/w_64_45# ALU_1b_1/AND_5/B 0.10fF
C3315 ALU_1b_3/AND_6/a_78_51# ALU_1b_3/AND_6/w_64_45# 0.09fF
C3316 ALU_1b_1/full_adder_0/w_448_45# vdd 0.12fF
C3317 gnd ALU_1b_2/AND_11/a_78_51# 0.07fF
C3318 ALU_1b_1/AND_15/A B3 0.28fF
C3319 ALU_1b_1/AND_16/a_78_51# gnd 0.07fF
C3320 gnd ALU_1b_2/AND_11/B 0.13fF
C3321 vdd ALU_1b_3/comparator_0/NOR_1/out 0.03fF
C3322 ALU_1b_1/AND_9/w_64_45# ALU_1b_1/AND_10/B 0.20fF
C3323 ALU_1b_2/AND_15/w_64_45# ALU_1b_2/NOR_1/B 0.06fF
C3324 ALU_1b_1/AND_2/w_64_45# ALU_1b_1/AND_2/B 0.06fF
C3325 ALU_1b_0/comparator_0/w_n195_n67# ALU_1b_0/comparator_0/NOR_3/out 0.11fF
C3326 vdd ALU_1b_2/comparator_0/AND_0/a_78_51# 0.06fF
C3327 ALU_1b_3/comparator_0/NOR_1/B ALU_1b_3/comparator_0/NOR_1/out 0.25fF
C3328 ALU_1b_2/AND_17/A ALU_1b_2/AND_17/a_78_51# 0.03fF
C3329 ALU_1b_1/NOT_4/in ALU_1b_1/NOR_2/B 0.15fF
C3330 ALU_1b_3/comparator_0/w_n195_n67# ALU_1b_3/comparator_0/NOR_3/B 0.06fF
C3331 ALU_1b_3/AND_8/out ALU_1b_3/C0 0.01fF
C3332 ALU_1b_0/decoder_0/AND_1/B ALU_1b_0/AND_2/B 0.17fF
C3333 ALU_1b_1/AND_2/out F2 0.01fF
C3334 vdd ALU_1b_3/NOR_3/B 0.33fF
C3335 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# ALU_1b_0/full_adder_0/NOR_0/B 0.12fF
C3336 ALU_1b_0/AND_17/w_64_45# ALU_1b_0/AND_17/a_78_51# 0.09fF
C3337 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# ALU_1b_1/AND_1/out 0.29fF
C3338 ALU_1b_2/comparator_0/AND_0/w_64_45# ALU_1b_2/comparator_0/AND_0/a_78_51# 0.09fF
C3339 ALU_1b_2/AND_6/out ALU_1b_2/comparator_0/AND_2/B 0.40fF
C3340 ALU_1b_3/AND_0/out ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# 0.13fF
C3341 S0 ALU_1b_3/decoder_0/AND_2/B 0.29fF
C3342 ALU_1b_0/AND_6/out ALU_1b_0/comparator_0/AND_1/a_78_51# 0.03fF
C3343 ALU_1b_0/comparator_0/AND_2/B ALU_1b_0/AND_9/out 0.29fF
C3344 ALU_1b_0/comparator_0/NOR_1/A gnd 0.17fF
C3345 ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out gnd 0.04fF
C3346 vdd ALU_1b_2/comparator_0/AND_3/w_64_45# 0.15fF
C3347 vdd ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_74# 0.02fF
C3348 ALU_1b_0/AND_9/out ALU_1b_0/AND_10/B 0.06fF
C3349 ALU_1b_2/AND_2/w_64_45# vdd 0.15fF
C3350 ALU_1b_3/AND_6/out ALU_1b_3/comparator_0/AND_1/w_64_45# 0.10fF
C3351 A0 ALU_1b_0/AND_12/w_64_45# 0.18fF
C3352 ALU_1b_3/AND_1/out ALU_1b_3/AND_16/A 0.11fF
C3353 ALU_1b_1/comparator_0/AND_1/w_64_45# ALU_1b_1/AND_9/out 0.39fF
C3354 ALU_1b_1/comparator_0/AND_2/B ALU_1b_1/comparator_0/AND_2/w_64_45# 0.06fF
C3355 gnd ALU_1b_2/comparator_0/AND_3/a_78_51# 0.07fF
C3356 ALU_1b_2/full_adder_0/w_448_45# ALU_1b_2/full_adder_0/NOR_0/out 0.11fF
C3357 ALU_1b_2/AND_1/a_78_51# ALU_1b_2/C0 0.03fF
C3358 ALU_1b_2/AND_1/out ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# 0.04fF
C3359 ALU_1b_0/AND_13/a_78_51# vdd 0.06fF
C3360 ALU_1b_2/full_adder_0/half_adder_1/A ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# 0.03fF
C3361 gnd ALU_1b_2/AND_5/B 0.48fF
C3362 ALU_1b_2/AND_2/out ALU_1b_2/full_adder_0/half_adder_1/A 0.11fF
C3363 ALU_1b_0/NOR_0/B ALU_1b_0/NOR_0/A 0.33fF
C3364 ALU_1b_0/AND_8/out gnd 0.23fF
C3365 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.09fF
C3366 ALU_1b_0/decoder_0/AND_1/B vdd 0.03fF
C3367 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# 0.22fF
C3368 vdd ALU_1b_2/NOR_2/w_n27_1# 0.24fF
C3369 ALU_1b_2/decoder_0/AND_3/a_78_51# ALU_1b_2/AND_12/w_64_45# 0.09fF
C3370 ALU_1b_3/AND_18/A ALU_1b_3/AND_18/a_78_51# 0.03fF
C3371 A0 ALU_1b_0/AND_5/B 0.01fF
C3372 ALU_1b_2/AND_3/out ALU_1b_2/AND_5/B 0.11fF
C3373 S0 ALU_1b_2/C0 0.22fF
C3374 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out ALU_1b_1/AND_5/out 0.20fF
C3375 ALU_1b_1/AND_9/w_64_45# vdd 0.42fF
C3376 ALU_1b_2/AND_0/out ALU_1b_2/C0 0.01fF
C3377 ALU_1b_0/AND_15/w_64_45# vdd 0.15fF
C3378 ALU_1b_0/AND_9/A vdd 1.07fF
C3379 ALU_1b_3/AND_2/a_78_51# B2 0.03fF
C3380 ALU_1b_2/AND_19/A ALU_1b_2/NOR_0/A 0.10fF
C3381 ALU_1b_1/full_adder_1/NOR_0/B ALU_1b_1/AND_3/out 0.10fF
C3382 ALU_1b_1/full_adder_1/NOR_0/A ALU_1b_1/NOT_1/in 0.23fF
C3383 ALU_1b_1/AND_10/a_78_51# gnd 0.07fF
C3384 vdd ALU_1b_3/decoder_0/AND_0/a_78_51# 0.06fF
C3385 ALU_1b_0/AND_15/a_78_51# gnd 0.07fF
C3386 ALU_1b_2/decoder_0/AND_2/a_78_51# ALU_1b_2/decoder_0/AND_2/B 0.19fF
C3387 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# vdd 0.06fF
C3388 ALU_1b_0/comparator_0/AND_2/a_78_51# ALU_1b_0/comparator_0/NOR_1/A 0.38fF
C3389 ALU_1b_2/AND_17/a_78_51# ALU_1b_2/AND_2/B 0.19fF
C3390 ALU_1b_1/AND_18/w_64_45# ALU_1b_1/NOR_3/A 0.03fF
C3391 ALU_1b_3/full_adder_1/half_adder_1/A ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# 0.00fF
C3392 ALU_1b_3/comparator_0/NOR_3/B ALU_1b_3/AND_8/out 0.02fF
C3393 ALU_1b_3/comparator_0/AND_2/w_64_45# ALU_1b_3/comparator_0/NOR_1/A 0.03fF
C3394 ALU_1b_1/comparator_0/NOR_3/B vdd 0.03fF
C3395 gnd ALU_1b_3/AND_3/out 0.11fF
C3396 ALU_1b_0/AND_1/w_64_45# ALU_1b_0/AND_2/B 0.06fF
C3397 ALU_1b_3/AND_10/a_78_51# ALU_1b_3/AND_9/A 0.05fF
C3398 ALU_1b_3/NOR_1/A ALU_1b_3/AND_11/B 0.03fF
C3399 ALU_1b_1/AND_0/out ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out 0.14fF
C3400 ALU_1b_0/AND_3/a_78_51# vdd 0.06fF
C3401 ALU_1b_1/decoder_0/AND_1/B S0 0.03fF
C3402 ALU_1b_1/comparator_0/NOR_3/out gnd 0.07fF
C3403 ALU_1b_2/comparator_0/AND_2/B ALU_1b_2/comparator_0/NOR_0/B 0.12fF
C3404 vdd ALU_1b_3/AND_6/out 0.20fF
C3405 ALU_1b_0/comparator_0/AND_1/a_78_51# ALU_1b_0/comparator_0/NOR_0/B 0.05fF
C3406 ALU_1b_0/comparator_0/AND_5/B ALU_1b_0/comparator_0/AND_5/a_78_51# 0.29fF
C3407 A1 ALU_1b_2/AND_9/A 0.31fF
C3408 ALU_1b_0/AND_14/w_64_45# ALU_1b_0/AND_13/a_78_51# 0.09fF
C3409 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_74# ALU_1b_3/NOT_1/in 0.03fF
C3410 ALU_1b_0/AND_7/a_78_51# ALU_1b_0/AND_9/A 0.05fF
C3411 vdd ALU_1b_2/NOR_0/B 0.20fF
C3412 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out gnd 0.04fF
C3413 ALU_1b_0/AND_1/a_78_51# ALU_1b_0/AND_2/B 0.19fF
C3414 gnd ALU_1b_3/decoder_0/AND_3/a_78_51# 0.07fF
C3415 ALU_1b_3/comparator_0/AND_5/B ALU_1b_3/comparator_0/AND_5/w_64_45# 0.06fF
C3416 ALU_1b_3/comparator_0/AND_1/w_64_45# ALU_1b_3/comparator_0/NOR_0/B 0.03fF
C3417 ALU_1b_0/NOR_1/A ALU_1b_0/NOR_2/A 0.12fF
C3418 ALU_1b_1/comparator_0/AND_2/w_64_45# vdd 0.15fF
C3419 ALU_1b_1/comparator_0/AND_5/w_64_45# ALU_1b_1/comparator_0/AND_5/a_78_51# 0.09fF
C3420 ALU_1b_1/comparator_0/AND_5/B ALU_1b_1/AND_7/out 0.61fF
C3421 ALU_1b_3/AND_7/w_64_45# ALU_1b_3/AND_9/A 0.39fF
C3422 ALU_1b_1/AND_13/a_78_51# ALU_1b_1/AND_15/A 0.05fF
C3423 ALU_1b_2/AND_1/out vdd 0.35fF
C3424 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# vdd 0.06fF
C3425 ALU_1b_1/AND_4/out ALU_1b_1/AND_5/out 0.11fF
C3426 ALU_1b_3/NOT_5/in ALU_1b_3/NOR_3/A 0.03fF
C3427 ALU_1b_1/AND_2/B ALU_1b_1/C0 0.28fF
C3428 ALU_1b_1/comparator_0/AND_2/a_78_51# gnd 0.07fF
C3429 ALU_1b_2/AND_3/w_64_45# ALU_1b_2/AND_5/B 0.06fF
C3430 ALU_1b_2/comparator_0/AND_5/w_64_45# ALU_1b_2/AND_7/out 0.30fF
C3431 ALU_1b_0/AND_17/A gnd 0.34fF
C3432 ALU_1b_0/AND_1/w_64_45# vdd 0.15fF
C3433 ALU_1b_0/comparator_0/AND_4/w_64_45# ALU_1b_0/AND_8/out 0.37fF
C3434 ALU_1b_2/AND_8/a_78_51# ALU_1b_2/AND_8/out 0.22fF
C3435 ALU_1b_0/AND_3/out Cin 0.01fF
C3436 ALU_1b_0/AND_14/B ALU_1b_0/AND_15/A 0.16fF
C3437 F0 ALU_1b_2/AND_5/B 0.01fF
C3438 ALU_1b_0/full_adder_1/w_448_45# vdd 0.12fF
C3439 ALU_1b_3/comparator_0/AND_2/B ALU_1b_3/comparator_0/w_n39_45# 0.03fF
C3440 ALU_1b_1/AND_15/w_64_45# ALU_1b_1/AND_15/A 0.06fF
C3441 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# vdd 0.06fF
C3442 gnd ALU_1b_2/NOR_3/A 0.23fF
C3443 ALU_1b_0/AND_1/a_78_51# vdd 0.06fF
C3444 ALU_1b_1/NOR_1/B ALU_1b_1/NOR_2/A 0.00fF
C3445 ALU_1b_2/full_adder_1/w_448_45# ALU_1b_2/full_adder_1/NOR_0/out 0.11fF
C3446 ALU_1b_0/AND_4/w_64_45# vdd 0.15fF
C3447 ALU_1b_2/AND_19/A ALU_1b_2/NOT_1/w_n36_43# 0.03fF
C3448 vdd ALU_1b_3/comparator_0/NOR_2/A 0.03fF
C3449 ALU_1b_0/full_adder_1/NOR_0/out gnd 0.07fF
C3450 ALU_1b_0/AND_4/a_78_51# gnd 0.07fF
C3451 gnd F1 0.38fF
C3452 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# ALU_1b_3/full_adder_0/half_adder_1/A 0.03fF
C3453 ALU_1b_3/NOR_0/B ALU_1b_3/NOT_2/in 0.15fF
C3454 ALU_1b_1/AND_14/B ALU_1b_1/AND_14/a_78_51# 0.19fF
C3455 ALU_1b_1/C0 ALU_1b_3/NOR_4/w_n27_1# 0.03fF
C3456 A3 ALU_1b_1/AND_6/w_64_45# 0.06fF
C3457 gnd ALU_1b_3/AND_17/A 0.34fF
C3458 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# 0.26fF
C3459 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# gnd 0.11fF
C3460 ALU_1b_0/AND_3/A vdd 0.03fF
C3461 vdd ALU_1b_3/comparator_0/NOR_0/B 0.09fF
C3462 ALU_1b_2/comparator_0/w_88_n67# ALU_1b_2/comparator_0/NOR_0/out 0.11fF
C3463 ALU_1b_1/AND_3/out ALU_1b_1/AND_4/a_78_51# 0.10fF
C3464 ALU_1b_0/comparator_0/NOR_0/out ALU_1b_0/comparator_0/NOR_1/B 0.05fF
C3465 vdd ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_74# 0.02fF
C3466 ALU_1b_3/AND_3/out ALU_1b_3/AND_4/out 0.98fF
C3467 ALU_1b_0/comparator_0/NOR_2/B ALU_1b_0/comparator_0/w_n195_n67# 0.19fF
C3468 vdd ALU_1b_2/comparator_0/w_n195_n67# 0.12fF
C3469 ALU_1b_3/comparator_0/NOR_0/B ALU_1b_3/comparator_0/NOR_1/B 0.01fF
C3470 gnd ALU_1b_3/comparator_0/NOR_0/out 0.07fF
C3471 ALU_1b_1/comparator_0/NOR_1/B ALU_1b_1/comparator_0/NOR_1/a_n14_7# 0.00fF
C3472 vdd ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_74# 0.02fF
C3473 ALU_1b_1/NOR_1/B vdd 0.20fF
C3474 ALU_1b_2/AND_2/w_64_45# B1 0.10fF
C3475 ALU_1b_3/full_adder_1/NOR_0/A ALU_1b_3/full_adder_1/half_adder_1/w_36_45# 0.03fF
C3476 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# vdd 0.06fF
C3477 ALU_1b_1/comparator_0/w_n195_n67# ALU_1b_1/comparator_0/NOR_3/A 0.06fF
C3478 ALU_1b_1/NOR_0/A ALU_1b_1/AND_5/B 0.01fF
C3479 ALU_1b_0/comparator_0/AND_1/w_64_45# vdd 0.14fF
C3480 ALU_1b_1/AND_13/a_78_51# B3 0.19fF
C3481 ALU_1b_1/comparator_0/NOR_2/B ALU_1b_1/AND_11/B 0.10fF
C3482 ALU_1b_0/full_adder_1/half_adder_1/A ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# 0.03fF
C3483 vdd ALU_1b_3/AND_16/a_78_51# 0.06fF
C3484 ALU_1b_1/AND_2/a_78_51# gnd 0.07fF
C3485 ALU_1b_0/comparator_0/AND_0/w_64_45# ALU_1b_0/comparator_0/AND_2/B 0.06fF
C3486 ALU_1b_0/comparator_0/AND_1/a_78_51# gnd 0.07fF
C3487 ALU_1b_2/AND_18/a_78_51# ALU_1b_2/AND_5/B 0.19fF
C3488 ALU_1b_3/AND_5/B Gnd 4.68fF
C3489 ALU_1b_3/NOT_3/in Gnd 0.42fF
C3490 ALU_1b_3/NOR_1/A Gnd 0.95fF
C3491 ALU_1b_3/NOR_2/w_n27_1# Gnd 2.18fF
C3492 F2 Gnd 1.52fF
C3493 ALU_1b_3/NOT_4/in Gnd 0.42fF
C3494 ALU_1b_3/NOT_2/in Gnd 0.42fF
C3495 ALU_1b_3/NOR_2/B Gnd 0.40fF
C3496 ALU_1b_3/AND_15/A Gnd 2.00fF
C3497 ALU_1b_3/decoder_0/AND_3/a_78_51# Gnd 0.42fF
C3498 ALU_1b_3/decoder_0/AND_2/a_78_51# Gnd 0.42fF
C3499 ALU_1b_3/decoder_0/AND_2/B Gnd 0.99fF
C3500 ALU_1b_3/AND_12/w_64_45# Gnd 3.63fF
C3501 ALU_1b_3/AND_9/A Gnd 3.01fF
C3502 ALU_1b_3/decoder_0/AND_1/a_78_51# Gnd 0.42fF
C3503 ALU_1b_3/decoder_0/AND_0/a_78_51# Gnd 0.42fF
C3504 ALU_1b_3/decoder_0/AND_1/B Gnd 1.73fF
C3505 ALU_1b_3/AND_6/w_64_45# Gnd 3.63fF
C3506 ALU_1b_3/NOR_2/A Gnd 0.06fF
C3507 ALU_1b_3/NOR_0/w_n27_1# Gnd 1.09fF
C3508 ALU_1b_3/AND_3/A Gnd 0.42fF
C3509 ALU_1b_3/NOT_1/w_n36_43# Gnd 0.48fF
C3510 ALU_1b_3/AND_10/B Gnd 1.14fF
C3511 ALU_1b_3/AND_11/B Gnd 1.00fF
C3512 ALU_1b_3/comparator_0/w_n39_45# Gnd 0.48fF
C3513 ALU_1b_3/comparator_0/w_n74_45# Gnd 0.48fF
C3514 ALU_1b_3/comparator_0/NOR_1/out Gnd 0.40fF
C3515 ALU_1b_3/comparator_0/NOR_1/B Gnd 1.06fF
C3516 ALU_1b_3/comparator_0/w_113_n67# Gnd 1.09fF
C3517 ALU_1b_3/comparator_0/NOR_0/out Gnd 0.40fF
C3518 ALU_1b_3/comparator_0/NOR_0/B Gnd 1.18fF
C3519 ALU_1b_3/comparator_0/w_88_n67# Gnd 1.09fF
C3520 ALU_1b_3/comparator_0/AND_4/a_78_51# Gnd 0.42fF
C3521 ALU_1b_3/AND_8/out Gnd 1.26fF
C3522 ALU_1b_3/AND_7/out Gnd 2.37fF
C3523 ALU_1b_3/comparator_0/AND_4/w_64_45# Gnd 1.05fF
C3524 ALU_1b_3/comparator_0/AND_5/a_78_51# Gnd 0.42fF
C3525 ALU_1b_3/comparator_0/AND_5/w_64_45# Gnd 1.05fF
C3526 ALU_1b_3/comparator_0/NOR_2/A Gnd 0.49fF
C3527 ALU_1b_3/comparator_0/AND_3/a_78_51# Gnd 0.42fF
C3528 ALU_1b_3/comparator_0/AND_5/B Gnd 0.66fF
C3529 ALU_1b_3/comparator_0/AND_3/w_64_45# Gnd 1.05fF
C3530 ALU_1b_3/comparator_0/NOR_1/A Gnd 0.97fF
C3531 ALU_1b_3/comparator_0/AND_2/a_78_51# Gnd 0.42fF
C3532 ALU_1b_3/comparator_0/AND_2/w_64_45# Gnd 1.05fF
C3533 ALU_1b_3/comparator_0/AND_1/a_78_51# Gnd 0.42fF
C3534 ALU_1b_3/AND_9/out Gnd 0.68fF
C3535 ALU_1b_3/comparator_0/AND_1/w_64_45# Gnd 1.05fF
C3536 ALU_1b_3/comparator_0/NOR_0/A Gnd 0.49fF
C3537 ALU_1b_3/comparator_0/AND_0/a_78_51# Gnd 0.42fF
C3538 ALU_1b_3/comparator_0/AND_2/B Gnd 0.66fF
C3539 ALU_1b_3/AND_6/out Gnd 1.12fF
C3540 ALU_1b_3/comparator_0/AND_0/w_64_45# Gnd 1.05fF
C3541 ALU_1b_3/comparator_0/NOR_3/out Gnd 0.11fF
C3542 ALU_1b_3/comparator_0/NOR_3/A Gnd 1.06fF
C3543 ALU_1b_3/comparator_0/w_n195_n67# Gnd 1.09fF
C3544 ALU_1b_3/comparator_0/NOR_2/out Gnd 0.40fF
C3545 ALU_1b_3/comparator_0/NOR_2/B Gnd 1.06fF
C3546 ALU_1b_3/comparator_0/w_n220_n67# Gnd 1.09fF
C3547 ALU_1b_3/NOR_3/A Gnd 0.53fF
C3548 ALU_1b_3/AND_18/a_78_51# Gnd 0.42fF
C3549 ALU_1b_3/AND_18/w_64_45# Gnd 1.05fF
C3550 ALU_1b_3/NOR_0/A Gnd 0.80fF
C3551 ALU_1b_3/AND_19/a_78_51# Gnd 0.42fF
C3552 ALU_1b_3/AND_19/A Gnd 0.62fF
C3553 ALU_1b_3/AND_19/w_64_45# Gnd 1.05fF
C3554 ALU_1b_3/NOR_3/B Gnd 0.66fF
C3555 ALU_1b_3/AND_17/a_78_51# Gnd 0.42fF
C3556 ALU_1b_3/AND_17/w_64_45# Gnd 1.05fF
C3557 ALU_1b_3/NOR_0/B Gnd 0.69fF
C3558 ALU_1b_3/AND_16/a_78_51# Gnd 0.42fF
C3559 ALU_1b_3/AND_16/w_64_45# Gnd 1.05fF
C3560 ALU_1b_3/NOR_1/B Gnd 0.58fF
C3561 ALU_1b_3/AND_15/a_78_51# Gnd 0.42fF
C3562 ALU_1b_3/AND_15/w_64_45# Gnd 1.05fF
C3563 ALU_1b_3/AND_15/B Gnd 0.79fF
C3564 ALU_1b_3/AND_14/a_78_51# Gnd 0.42fF
C3565 ALU_1b_3/AND_14/B Gnd 0.93fF
C3566 ALU_1b_3/AND_14/A Gnd 0.42fF
C3567 ALU_1b_3/AND_9/a_78_51# Gnd 0.42fF
C3568 ALU_1b_3/AND_13/a_78_51# Gnd 0.42fF
C3569 ALU_1b_3/AND_14/w_64_45# Gnd 2.10fF
C3570 ALU_1b_3/AND_8/a_78_51# Gnd 0.42fF
C3571 ALU_1b_3/AND_8/w_64_45# Gnd 1.05fF
C3572 ALU_1b_3/AND_12/a_78_51# Gnd 0.42fF
C3573 ALU_1b_3/AND_7/a_78_51# Gnd 0.42fF
C3574 ALU_1b_3/AND_7/w_64_45# Gnd 1.05fF
C3575 ALU_1b_3/AND_6/a_78_51# Gnd 0.42fF
C3576 ALU_1b_3/AND_11/a_78_51# Gnd 0.42fF
C3577 ALU_1b_3/AND_10/a_78_51# Gnd 0.42fF
C3578 ALU_1b_3/AND_9/w_64_45# Gnd 3.15fF
C3579 ALU_1b_3/AND_4/a_78_51# Gnd 0.42fF
C3580 ALU_1b_3/AND_4/w_64_45# Gnd 1.05fF
C3581 ALU_1b_3/AND_5/a_78_51# Gnd 0.42fF
C3582 ALU_1b_3/AND_5/w_64_45# Gnd 1.05fF
C3583 ALU_1b_3/AND_3/a_78_51# Gnd 0.42fF
C3584 ALU_1b_3/AND_3/w_64_45# Gnd 1.53fF
C3585 ALU_1b_3/AND_2/a_78_51# Gnd 0.42fF
C3586 ALU_1b_3/AND_2/w_64_45# Gnd 1.05fF
C3587 ALU_1b_3/AND_18/A Gnd 0.73fF
C3588 ALU_1b_3/full_adder_1/NOR_0/out Gnd 0.39fF
C3589 ALU_1b_3/full_adder_1/w_448_45# Gnd 1.07fF
C3590 ALU_1b_3/full_adder_1/NOR_0/B Gnd 0.74fF
C3591 ALU_1b_3/AND_4/out Gnd 1.58fF
C3592 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3593 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3594 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3595 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3596 ALU_1b_3/AND_3/out Gnd 2.67fF
C3597 ALU_1b_3/full_adder_1/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3598 ALU_1b_3/full_adder_1/half_adder_0/NAND_0/out Gnd 0.43fF
C3599 ALU_1b_3/full_adder_1/half_adder_0/w_36_45# Gnd 1.11fF
C3600 ALU_1b_3/full_adder_1/NOR_0/A Gnd 0.64fF
C3601 ALU_1b_3/AND_5/out Gnd 2.18fF
C3602 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3603 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3604 ALU_1b_3/NOT_1/in Gnd 1.41fF
C3605 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3606 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3607 ALU_1b_3/full_adder_1/half_adder_1/A Gnd 2.66fF
C3608 ALU_1b_3/full_adder_1/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3609 ALU_1b_3/full_adder_1/half_adder_1/NAND_0/out Gnd 0.43fF
C3610 ALU_1b_3/full_adder_1/half_adder_1/w_36_45# Gnd 1.11fF
C3611 ALU_1b_3/AND_1/a_78_51# Gnd 0.42fF
C3612 ALU_1b_3/AND_1/w_64_45# Gnd 1.05fF
C3613 ALU_1b_3/AND_17/A Gnd 0.81fF
C3614 ALU_1b_3/full_adder_0/NOR_0/out Gnd 0.39fF
C3615 ALU_1b_3/full_adder_0/w_448_45# Gnd 1.07fF
C3616 ALU_1b_3/full_adder_0/NOR_0/B Gnd 0.74fF
C3617 ALU_1b_3/AND_2/out Gnd 1.53fF
C3618 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3619 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3620 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3621 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3622 ALU_1b_3/AND_0/out Gnd 3.03fF
C3623 ALU_1b_3/full_adder_0/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3624 ALU_1b_3/full_adder_0/half_adder_0/NAND_0/out Gnd 0.43fF
C3625 ALU_1b_3/full_adder_0/half_adder_0/w_36_45# Gnd 1.11fF
C3626 ALU_1b_3/full_adder_0/NOR_0/A Gnd 0.64fF
C3627 ALU_1b_3/AND_1/out Gnd 2.07fF
C3628 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3629 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3630 ALU_1b_3/AND_16/A Gnd 1.26fF
C3631 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3632 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3633 ALU_1b_3/full_adder_0/half_adder_1/A Gnd 2.66fF
C3634 ALU_1b_3/full_adder_0/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3635 ALU_1b_3/full_adder_0/half_adder_1/NAND_0/out Gnd 0.43fF
C3636 ALU_1b_3/full_adder_0/half_adder_1/w_36_45# Gnd 1.11fF
C3637 ALU_1b_3/AND_0/a_78_51# Gnd 0.42fF
C3638 ALU_1b_3/AND_0/w_64_45# Gnd 1.05fF
C3639 ALU_1b_3/NOT_6/in Gnd 0.42fF
C3640 ALU_1b_3/NOR_4/B Gnd 0.40fF
C3641 ALU_1b_3/NOR_4/A Gnd 0.82fF
C3642 ALU_1b_3/NOT_5/in Gnd 0.42fF
C3643 ALU_1b_3/NOR_4/w_n27_1# Gnd 2.18fF
C3644 ALU_1b_2/AND_5/B Gnd 4.68fF
C3645 ALU_1b_2/NOT_3/in Gnd 0.42fF
C3646 ALU_1b_2/NOR_1/A Gnd 0.95fF
C3647 ALU_1b_2/NOR_2/w_n27_1# Gnd 2.18fF
C3648 ALU_1b_2/NOT_4/in Gnd 0.42fF
C3649 ALU_1b_2/NOT_2/in Gnd 0.42fF
C3650 ALU_1b_2/NOR_2/B Gnd 0.40fF
C3651 ALU_1b_2/AND_15/A Gnd 2.00fF
C3652 ALU_1b_2/decoder_0/AND_3/a_78_51# Gnd 0.42fF
C3653 ALU_1b_2/decoder_0/AND_2/a_78_51# Gnd 0.42fF
C3654 ALU_1b_2/decoder_0/AND_2/B Gnd 0.99fF
C3655 ALU_1b_2/AND_12/w_64_45# Gnd 3.63fF
C3656 ALU_1b_2/AND_9/A Gnd 3.01fF
C3657 ALU_1b_2/decoder_0/AND_1/a_78_51# Gnd 0.42fF
C3658 ALU_1b_2/decoder_0/AND_0/a_78_51# Gnd 0.42fF
C3659 ALU_1b_2/decoder_0/AND_1/B Gnd 1.73fF
C3660 ALU_1b_2/AND_6/w_64_45# Gnd 3.63fF
C3661 ALU_1b_2/NOR_2/A Gnd 0.06fF
C3662 ALU_1b_2/NOR_0/w_n27_1# Gnd 1.09fF
C3663 ALU_1b_2/AND_3/A Gnd 0.42fF
C3664 ALU_1b_2/NOT_1/w_n36_43# Gnd 0.48fF
C3665 ALU_1b_2/AND_10/B Gnd 1.14fF
C3666 ALU_1b_2/AND_11/B Gnd 1.00fF
C3667 ALU_1b_2/comparator_0/w_n39_45# Gnd 0.48fF
C3668 ALU_1b_2/comparator_0/w_n74_45# Gnd 0.48fF
C3669 ALU_1b_2/comparator_0/NOR_1/out Gnd 0.40fF
C3670 ALU_1b_2/comparator_0/NOR_1/B Gnd 1.06fF
C3671 ALU_1b_2/comparator_0/w_113_n67# Gnd 1.09fF
C3672 ALU_1b_2/comparator_0/NOR_0/out Gnd 0.40fF
C3673 ALU_1b_2/comparator_0/NOR_0/B Gnd 1.18fF
C3674 ALU_1b_2/comparator_0/w_88_n67# Gnd 1.09fF
C3675 ALU_1b_2/comparator_0/AND_4/a_78_51# Gnd 0.42fF
C3676 ALU_1b_2/AND_8/out Gnd 1.26fF
C3677 ALU_1b_2/AND_7/out Gnd 2.37fF
C3678 ALU_1b_2/comparator_0/AND_4/w_64_45# Gnd 1.05fF
C3679 ALU_1b_2/comparator_0/AND_5/a_78_51# Gnd 0.42fF
C3680 ALU_1b_2/comparator_0/AND_5/w_64_45# Gnd 1.05fF
C3681 ALU_1b_2/comparator_0/NOR_2/A Gnd 0.49fF
C3682 ALU_1b_2/comparator_0/AND_3/a_78_51# Gnd 0.42fF
C3683 ALU_1b_2/comparator_0/AND_5/B Gnd 0.66fF
C3684 ALU_1b_2/comparator_0/AND_3/w_64_45# Gnd 1.05fF
C3685 ALU_1b_2/comparator_0/NOR_1/A Gnd 0.97fF
C3686 ALU_1b_2/comparator_0/AND_2/a_78_51# Gnd 0.42fF
C3687 ALU_1b_2/comparator_0/AND_2/w_64_45# Gnd 1.05fF
C3688 ALU_1b_2/comparator_0/AND_1/a_78_51# Gnd 0.42fF
C3689 ALU_1b_2/AND_9/out Gnd 0.68fF
C3690 ALU_1b_2/comparator_0/AND_1/w_64_45# Gnd 1.05fF
C3691 ALU_1b_2/comparator_0/NOR_0/A Gnd 0.49fF
C3692 ALU_1b_2/comparator_0/AND_0/a_78_51# Gnd 0.42fF
C3693 ALU_1b_2/comparator_0/AND_2/B Gnd 0.66fF
C3694 ALU_1b_2/AND_6/out Gnd 1.12fF
C3695 ALU_1b_2/comparator_0/AND_0/w_64_45# Gnd 1.05fF
C3696 ALU_1b_2/comparator_0/NOR_3/out Gnd 0.11fF
C3697 ALU_1b_2/comparator_0/NOR_3/A Gnd 1.06fF
C3698 ALU_1b_2/comparator_0/w_n195_n67# Gnd 1.09fF
C3699 ALU_1b_2/comparator_0/NOR_2/out Gnd 0.40fF
C3700 ALU_1b_2/comparator_0/NOR_2/B Gnd 1.06fF
C3701 ALU_1b_2/comparator_0/w_n220_n67# Gnd 1.09fF
C3702 ALU_1b_2/NOR_3/A Gnd 0.53fF
C3703 ALU_1b_2/AND_18/a_78_51# Gnd 0.42fF
C3704 ALU_1b_2/AND_18/w_64_45# Gnd 1.05fF
C3705 ALU_1b_2/NOR_0/A Gnd 0.80fF
C3706 ALU_1b_2/AND_19/a_78_51# Gnd 0.42fF
C3707 ALU_1b_2/AND_19/A Gnd 0.62fF
C3708 ALU_1b_2/AND_19/w_64_45# Gnd 1.05fF
C3709 ALU_1b_2/NOR_3/B Gnd 0.66fF
C3710 ALU_1b_2/AND_17/a_78_51# Gnd 0.42fF
C3711 ALU_1b_2/AND_17/w_64_45# Gnd 1.05fF
C3712 ALU_1b_2/NOR_0/B Gnd 0.69fF
C3713 ALU_1b_2/AND_16/a_78_51# Gnd 0.42fF
C3714 ALU_1b_2/AND_16/w_64_45# Gnd 1.05fF
C3715 ALU_1b_2/NOR_1/B Gnd 0.58fF
C3716 ALU_1b_2/AND_15/a_78_51# Gnd 0.42fF
C3717 ALU_1b_2/AND_15/w_64_45# Gnd 1.05fF
C3718 ALU_1b_2/AND_15/B Gnd 0.79fF
C3719 ALU_1b_2/AND_14/a_78_51# Gnd 0.42fF
C3720 ALU_1b_2/AND_14/B Gnd 0.93fF
C3721 ALU_1b_2/AND_14/A Gnd 0.42fF
C3722 ALU_1b_2/AND_9/a_78_51# Gnd 0.42fF
C3723 F0 Gnd 1.57fF
C3724 ALU_1b_2/AND_13/a_78_51# Gnd 0.42fF
C3725 ALU_1b_2/AND_14/w_64_45# Gnd 2.10fF
C3726 ALU_1b_2/AND_8/a_78_51# Gnd 0.42fF
C3727 ALU_1b_2/AND_8/w_64_45# Gnd 1.05fF
C3728 ALU_1b_2/AND_12/a_78_51# Gnd 0.42fF
C3729 ALU_1b_2/AND_7/a_78_51# Gnd 0.42fF
C3730 ALU_1b_2/AND_7/w_64_45# Gnd 1.05fF
C3731 ALU_1b_2/AND_6/a_78_51# Gnd 0.42fF
C3732 ALU_1b_2/AND_11/a_78_51# Gnd 0.42fF
C3733 ALU_1b_2/AND_10/a_78_51# Gnd 0.42fF
C3734 ALU_1b_2/AND_9/w_64_45# Gnd 3.15fF
C3735 ALU_1b_2/AND_4/a_78_51# Gnd 0.42fF
C3736 ALU_1b_2/AND_4/w_64_45# Gnd 1.05fF
C3737 ALU_1b_2/AND_5/a_78_51# Gnd 0.42fF
C3738 ALU_1b_2/AND_5/w_64_45# Gnd 1.05fF
C3739 ALU_1b_2/AND_3/a_78_51# Gnd 0.42fF
C3740 ALU_1b_2/AND_3/w_64_45# Gnd 1.53fF
C3741 ALU_1b_2/AND_2/a_78_51# Gnd 0.42fF
C3742 ALU_1b_2/AND_2/w_64_45# Gnd 1.05fF
C3743 ALU_1b_2/AND_18/A Gnd 0.73fF
C3744 ALU_1b_2/full_adder_1/NOR_0/out Gnd 0.39fF
C3745 ALU_1b_2/full_adder_1/w_448_45# Gnd 1.07fF
C3746 ALU_1b_2/full_adder_1/NOR_0/B Gnd 0.74fF
C3747 ALU_1b_2/AND_4/out Gnd 1.58fF
C3748 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3749 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3750 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3751 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3752 ALU_1b_2/AND_3/out Gnd 2.67fF
C3753 ALU_1b_2/full_adder_1/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3754 ALU_1b_2/full_adder_1/half_adder_0/NAND_0/out Gnd 0.43fF
C3755 ALU_1b_2/full_adder_1/half_adder_0/w_36_45# Gnd 1.11fF
C3756 ALU_1b_2/full_adder_1/NOR_0/A Gnd 0.64fF
C3757 ALU_1b_2/AND_5/out Gnd 2.18fF
C3758 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3759 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3760 ALU_1b_2/NOT_1/in Gnd 1.41fF
C3761 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3762 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3763 ALU_1b_2/full_adder_1/half_adder_1/A Gnd 2.66fF
C3764 ALU_1b_2/full_adder_1/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3765 ALU_1b_2/full_adder_1/half_adder_1/NAND_0/out Gnd 0.43fF
C3766 ALU_1b_2/full_adder_1/half_adder_1/w_36_45# Gnd 1.11fF
C3767 ALU_1b_2/AND_1/a_78_51# Gnd 0.42fF
C3768 ALU_1b_2/AND_1/w_64_45# Gnd 1.05fF
C3769 ALU_1b_2/AND_17/A Gnd 0.81fF
C3770 ALU_1b_2/full_adder_0/NOR_0/out Gnd 0.39fF
C3771 ALU_1b_2/full_adder_0/w_448_45# Gnd 1.07fF
C3772 ALU_1b_2/full_adder_0/NOR_0/B Gnd 0.74fF
C3773 ALU_1b_2/AND_2/out Gnd 1.53fF
C3774 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3775 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3776 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3777 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3778 ALU_1b_2/AND_0/out Gnd 3.03fF
C3779 ALU_1b_2/full_adder_0/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3780 ALU_1b_2/full_adder_0/half_adder_0/NAND_0/out Gnd 0.43fF
C3781 ALU_1b_2/full_adder_0/half_adder_0/w_36_45# Gnd 1.11fF
C3782 ALU_1b_2/full_adder_0/NOR_0/A Gnd 0.64fF
C3783 ALU_1b_2/AND_1/out Gnd 2.07fF
C3784 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3785 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3786 ALU_1b_2/AND_16/A Gnd 1.26fF
C3787 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3788 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3789 ALU_1b_2/full_adder_0/half_adder_1/A Gnd 2.66fF
C3790 ALU_1b_2/full_adder_0/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3791 ALU_1b_2/full_adder_0/half_adder_1/NAND_0/out Gnd 0.43fF
C3792 ALU_1b_2/full_adder_0/half_adder_1/w_36_45# Gnd 1.11fF
C3793 ALU_1b_2/AND_0/a_78_51# Gnd 0.42fF
C3794 ALU_1b_2/AND_0/w_64_45# Gnd 1.05fF
C3795 ALU_1b_2/NOT_6/in Gnd 0.42fF
C3796 ALU_1b_2/NOR_4/B Gnd 0.40fF
C3797 ALU_1b_2/NOR_4/A Gnd 0.82fF
C3798 ALU_1b_2/NOT_5/in Gnd 0.42fF
C3799 ALU_1b_2/NOR_4/w_n27_1# Gnd 2.18fF
C3800 gnd Gnd 86.94fF
C3801 ALU_1b_1/AND_5/B Gnd 4.68fF
C3802 ALU_1b_1/NOT_3/in Gnd 0.42fF
C3803 ALU_1b_1/NOR_1/A Gnd 0.95fF
C3804 ALU_1b_1/NOR_2/w_n27_1# Gnd 2.18fF
C3805 F3 Gnd 0.56fF
C3806 ALU_1b_1/NOT_4/in Gnd 0.42fF
C3807 ALU_1b_1/NOT_2/in Gnd 0.42fF
C3808 ALU_1b_1/NOR_2/B Gnd 0.40fF
C3809 ALU_1b_1/AND_15/A Gnd 2.00fF
C3810 ALU_1b_1/decoder_0/AND_3/a_78_51# Gnd 0.42fF
C3811 ALU_1b_1/decoder_0/AND_2/a_78_51# Gnd 0.42fF
C3812 ALU_1b_1/decoder_0/AND_2/B Gnd 0.99fF
C3813 ALU_1b_1/AND_12/w_64_45# Gnd 3.63fF
C3814 ALU_1b_1/AND_9/A Gnd 3.01fF
C3815 ALU_1b_1/decoder_0/AND_1/a_78_51# Gnd 0.42fF
C3816 ALU_1b_1/decoder_0/AND_0/a_78_51# Gnd 0.42fF
C3817 ALU_1b_1/decoder_0/AND_1/B Gnd 1.73fF
C3818 ALU_1b_1/AND_6/w_64_45# Gnd 3.63fF
C3819 ALU_1b_1/NOR_2/A Gnd 0.06fF
C3820 ALU_1b_1/NOR_0/w_n27_1# Gnd 1.09fF
C3821 ALU_1b_1/AND_3/A Gnd 0.42fF
C3822 ALU_1b_1/NOT_1/w_n36_43# Gnd 0.48fF
C3823 ALU_1b_1/AND_10/B Gnd 1.14fF
C3824 ALU_1b_1/AND_11/B Gnd 1.00fF
C3825 ALU_1b_1/comparator_0/w_n39_45# Gnd 0.48fF
C3826 ALU_1b_1/comparator_0/w_n74_45# Gnd 0.48fF
C3827 ALU_1b_1/comparator_0/NOR_1/out Gnd 0.40fF
C3828 ALU_1b_1/comparator_0/NOR_1/B Gnd 1.06fF
C3829 ALU_1b_1/comparator_0/w_113_n67# Gnd 1.09fF
C3830 ALU_1b_1/comparator_0/NOR_0/out Gnd 0.40fF
C3831 vdd Gnd 31.71fF
C3832 ALU_1b_1/comparator_0/NOR_0/B Gnd 1.18fF
C3833 ALU_1b_1/comparator_0/w_88_n67# Gnd 1.09fF
C3834 ALU_1b_1/comparator_0/AND_4/a_78_51# Gnd 0.42fF
C3835 ALU_1b_1/AND_8/out Gnd 1.26fF
C3836 ALU_1b_1/AND_7/out Gnd 2.37fF
C3837 ALU_1b_1/comparator_0/AND_4/w_64_45# Gnd 1.05fF
C3838 ALU_1b_1/comparator_0/AND_5/a_78_51# Gnd 0.42fF
C3839 ALU_1b_1/comparator_0/AND_5/w_64_45# Gnd 1.05fF
C3840 ALU_1b_1/comparator_0/NOR_2/A Gnd 0.49fF
C3841 ALU_1b_1/comparator_0/AND_3/a_78_51# Gnd 0.42fF
C3842 ALU_1b_1/comparator_0/AND_5/B Gnd 0.66fF
C3843 ALU_1b_1/comparator_0/AND_3/w_64_45# Gnd 1.05fF
C3844 ALU_1b_1/comparator_0/NOR_1/A Gnd 0.97fF
C3845 ALU_1b_1/comparator_0/AND_2/a_78_51# Gnd 0.42fF
C3846 ALU_1b_1/comparator_0/AND_2/w_64_45# Gnd 1.05fF
C3847 ALU_1b_1/comparator_0/AND_1/a_78_51# Gnd 0.42fF
C3848 ALU_1b_1/AND_9/out Gnd 0.68fF
C3849 ALU_1b_1/comparator_0/AND_1/w_64_45# Gnd 1.05fF
C3850 ALU_1b_1/comparator_0/NOR_0/A Gnd 0.49fF
C3851 ALU_1b_1/comparator_0/AND_0/a_78_51# Gnd 0.42fF
C3852 ALU_1b_1/comparator_0/AND_2/B Gnd 0.66fF
C3853 ALU_1b_1/AND_6/out Gnd 1.12fF
C3854 ALU_1b_1/comparator_0/AND_0/w_64_45# Gnd 1.05fF
C3855 ALU_1b_1/comparator_0/NOR_3/out Gnd 0.11fF
C3856 ALU_1b_1/comparator_0/NOR_3/A Gnd 1.06fF
C3857 ALU_1b_1/comparator_0/w_n195_n67# Gnd 1.09fF
C3858 ALU_1b_1/comparator_0/NOR_2/out Gnd 0.40fF
C3859 ALU_1b_1/comparator_0/NOR_2/B Gnd 1.06fF
C3860 ALU_1b_1/comparator_0/w_n220_n67# Gnd 1.09fF
C3861 ALU_1b_1/NOR_3/A Gnd 0.53fF
C3862 ALU_1b_1/AND_18/a_78_51# Gnd 0.42fF
C3863 ALU_1b_1/AND_18/w_64_45# Gnd 1.05fF
C3864 ALU_1b_1/NOR_0/A Gnd 0.80fF
C3865 ALU_1b_1/AND_19/a_78_51# Gnd 0.42fF
C3866 ALU_1b_1/AND_19/A Gnd 0.62fF
C3867 ALU_1b_1/AND_19/w_64_45# Gnd 1.05fF
C3868 ALU_1b_1/NOR_3/B Gnd 0.66fF
C3869 ALU_1b_1/AND_17/a_78_51# Gnd 0.42fF
C3870 ALU_1b_1/AND_17/w_64_45# Gnd 1.05fF
C3871 ALU_1b_1/NOR_0/B Gnd 0.69fF
C3872 ALU_1b_1/AND_16/a_78_51# Gnd 0.42fF
C3873 ALU_1b_1/AND_16/w_64_45# Gnd 1.05fF
C3874 ALU_1b_1/NOR_1/B Gnd 0.58fF
C3875 ALU_1b_1/AND_15/a_78_51# Gnd 0.42fF
C3876 ALU_1b_1/AND_15/w_64_45# Gnd 1.05fF
C3877 ALU_1b_1/AND_15/B Gnd 0.79fF
C3878 ALU_1b_1/AND_14/a_78_51# Gnd 0.42fF
C3879 ALU_1b_1/AND_14/B Gnd 0.93fF
C3880 ALU_1b_1/AND_14/A Gnd 0.42fF
C3881 ALU_1b_1/AND_9/a_78_51# Gnd 0.42fF
C3882 ALU_1b_1/AND_13/a_78_51# Gnd 0.42fF
C3883 ALU_1b_1/AND_14/w_64_45# Gnd 2.10fF
C3884 ALU_1b_1/AND_8/a_78_51# Gnd 0.42fF
C3885 ALU_1b_1/AND_8/w_64_45# Gnd 1.05fF
C3886 ALU_1b_1/AND_12/a_78_51# Gnd 0.42fF
C3887 ALU_1b_1/AND_7/a_78_51# Gnd 0.42fF
C3888 ALU_1b_1/AND_7/w_64_45# Gnd 1.05fF
C3889 ALU_1b_1/AND_6/a_78_51# Gnd 0.42fF
C3890 ALU_1b_1/AND_11/a_78_51# Gnd 0.42fF
C3891 ALU_1b_1/AND_10/a_78_51# Gnd 0.42fF
C3892 ALU_1b_1/AND_9/w_64_45# Gnd 3.15fF
C3893 ALU_1b_1/AND_4/a_78_51# Gnd 0.42fF
C3894 ALU_1b_1/AND_4/w_64_45# Gnd 1.05fF
C3895 ALU_1b_1/AND_5/a_78_51# Gnd 0.42fF
C3896 ALU_1b_1/AND_5/w_64_45# Gnd 1.05fF
C3897 ALU_1b_1/AND_3/a_78_51# Gnd 0.42fF
C3898 ALU_1b_1/AND_3/w_64_45# Gnd 1.53fF
C3899 ALU_1b_1/AND_2/a_78_51# Gnd 0.42fF
C3900 ALU_1b_1/AND_2/w_64_45# Gnd 1.05fF
C3901 ALU_1b_1/AND_18/A Gnd 0.73fF
C3902 ALU_1b_1/full_adder_1/NOR_0/out Gnd 0.39fF
C3903 ALU_1b_1/full_adder_1/w_448_45# Gnd 1.07fF
C3904 ALU_1b_1/full_adder_1/NOR_0/B Gnd 0.74fF
C3905 ALU_1b_1/AND_4/out Gnd 1.58fF
C3906 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3907 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3908 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3909 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3910 ALU_1b_1/AND_3/out Gnd 2.67fF
C3911 ALU_1b_1/full_adder_1/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3912 ALU_1b_1/full_adder_1/half_adder_0/NAND_0/out Gnd 0.43fF
C3913 ALU_1b_1/full_adder_1/half_adder_0/w_36_45# Gnd 1.11fF
C3914 ALU_1b_1/full_adder_1/NOR_0/A Gnd 0.64fF
C3915 ALU_1b_1/AND_5/out Gnd 2.18fF
C3916 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3917 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3918 ALU_1b_1/NOT_1/in Gnd 1.41fF
C3919 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3920 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3921 ALU_1b_1/full_adder_1/half_adder_1/A Gnd 2.66fF
C3922 ALU_1b_1/full_adder_1/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3923 ALU_1b_1/full_adder_1/half_adder_1/NAND_0/out Gnd 0.43fF
C3924 ALU_1b_1/full_adder_1/half_adder_1/w_36_45# Gnd 1.11fF
C3925 ALU_1b_1/AND_1/a_78_51# Gnd 0.42fF
C3926 ALU_1b_1/AND_1/w_64_45# Gnd 1.05fF
C3927 ALU_1b_1/AND_17/A Gnd 0.81fF
C3928 ALU_1b_1/full_adder_0/NOR_0/out Gnd 0.39fF
C3929 ALU_1b_1/full_adder_0/w_448_45# Gnd 1.07fF
C3930 ALU_1b_1/full_adder_0/NOR_0/B Gnd 0.74fF
C3931 ALU_1b_1/AND_2/out Gnd 1.53fF
C3932 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C3933 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C3934 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C3935 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C3936 ALU_1b_1/AND_0/out Gnd 3.03fF
C3937 ALU_1b_1/full_adder_0/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C3938 ALU_1b_1/full_adder_0/half_adder_0/NAND_0/out Gnd 0.43fF
C3939 ALU_1b_1/full_adder_0/half_adder_0/w_36_45# Gnd 1.11fF
C3940 ALU_1b_1/full_adder_0/NOR_0/A Gnd 0.64fF
C3941 ALU_1b_1/AND_1/out Gnd 2.07fF
C3942 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C3943 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C3944 ALU_1b_1/AND_16/A Gnd 1.26fF
C3945 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C3946 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C3947 ALU_1b_1/full_adder_0/half_adder_1/A Gnd 2.66fF
C3948 ALU_1b_1/full_adder_0/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C3949 ALU_1b_1/full_adder_0/half_adder_1/NAND_0/out Gnd 0.43fF
C3950 ALU_1b_1/full_adder_0/half_adder_1/w_36_45# Gnd 1.11fF
C3951 ALU_1b_1/AND_0/a_78_51# Gnd 0.42fF
C3952 ALU_1b_1/AND_0/w_64_45# Gnd 1.05fF
C3953 ALU_1b_1/NOT_6/in Gnd 0.42fF
C3954 ALU_1b_1/NOR_4/B Gnd 0.40fF
C3955 ALU_1b_1/NOR_4/A Gnd 0.82fF
C3956 ALU_1b_1/NOT_5/in Gnd 0.42fF
C3957 ALU_1b_1/NOR_4/w_n27_1# Gnd 2.18fF
C3958 ALU_1b_0/AND_5/B Gnd 4.68fF
C3959 ALU_1b_0/NOT_3/in Gnd 0.42fF
C3960 ALU_1b_0/NOR_1/A Gnd 0.95fF
C3961 ALU_1b_0/NOR_2/w_n27_1# Gnd 2.18fF
C3962 ALU_1b_0/NOT_4/in Gnd 0.42fF
C3963 ALU_1b_0/NOT_2/in Gnd 0.42fF
C3964 ALU_1b_0/NOR_2/B Gnd 0.40fF
C3965 ALU_1b_0/AND_15/A Gnd 2.00fF
C3966 ALU_1b_0/decoder_0/AND_3/a_78_51# Gnd 0.42fF
C3967 ALU_1b_0/decoder_0/AND_2/a_78_51# Gnd 0.42fF
C3968 ALU_1b_0/decoder_0/AND_2/B Gnd 0.99fF
C3969 ALU_1b_0/AND_12/w_64_45# Gnd 3.63fF
C3970 ALU_1b_0/AND_9/A Gnd 3.01fF
C3971 ALU_1b_0/decoder_0/AND_1/a_78_51# Gnd 0.42fF
C3972 ALU_1b_0/decoder_0/AND_0/a_78_51# Gnd 0.42fF
C3973 ALU_1b_0/decoder_0/AND_1/B Gnd 1.73fF
C3974 ALU_1b_0/AND_6/w_64_45# Gnd 3.63fF
C3975 ALU_1b_0/NOR_2/A Gnd 0.06fF
C3976 ALU_1b_0/NOR_0/w_n27_1# Gnd 1.09fF
C3977 ALU_1b_0/AND_3/A Gnd 0.42fF
C3978 ALU_1b_0/NOT_1/w_n36_43# Gnd 0.48fF
C3979 ALU_1b_0/AND_10/B Gnd 1.14fF
C3980 ALU_1b_0/AND_11/B Gnd 1.00fF
C3981 ALU_1b_0/comparator_0/w_n39_45# Gnd 0.48fF
C3982 ALU_1b_0/comparator_0/w_n74_45# Gnd 0.48fF
C3983 ALU_1b_0/comparator_0/NOR_1/out Gnd 0.40fF
C3984 ALU_1b_0/comparator_0/NOR_1/B Gnd 1.06fF
C3985 ALU_1b_0/comparator_0/w_113_n67# Gnd 1.09fF
C3986 ALU_1b_0/comparator_0/NOR_0/out Gnd 0.40fF
C3987 ALU_1b_0/comparator_0/NOR_0/B Gnd 1.18fF
C3988 ALU_1b_0/comparator_0/w_88_n67# Gnd 1.09fF
C3989 ALU_1b_0/comparator_0/AND_4/a_78_51# Gnd 0.42fF
C3990 ALU_1b_0/AND_8/out Gnd 1.26fF
C3991 ALU_1b_0/AND_7/out Gnd 2.37fF
C3992 ALU_1b_0/comparator_0/AND_4/w_64_45# Gnd 1.05fF
C3993 ALU_1b_0/comparator_0/AND_5/a_78_51# Gnd 0.42fF
C3994 ALU_1b_0/comparator_0/AND_5/w_64_45# Gnd 1.05fF
C3995 ALU_1b_0/comparator_0/NOR_2/A Gnd 0.49fF
C3996 ALU_1b_0/comparator_0/AND_3/a_78_51# Gnd 0.42fF
C3997 ALU_1b_0/comparator_0/AND_5/B Gnd 0.66fF
C3998 ALU_1b_0/comparator_0/AND_3/w_64_45# Gnd 1.05fF
C3999 ALU_1b_0/comparator_0/NOR_1/A Gnd 0.97fF
C4000 ALU_1b_0/comparator_0/AND_2/a_78_51# Gnd 0.42fF
C4001 ALU_1b_0/comparator_0/AND_2/w_64_45# Gnd 1.05fF
C4002 ALU_1b_0/comparator_0/AND_1/a_78_51# Gnd 0.42fF
C4003 ALU_1b_0/AND_9/out Gnd 0.68fF
C4004 ALU_1b_0/comparator_0/AND_1/w_64_45# Gnd 1.05fF
C4005 ALU_1b_0/comparator_0/NOR_0/A Gnd 0.49fF
C4006 ALU_1b_0/comparator_0/AND_0/a_78_51# Gnd 0.42fF
C4007 ALU_1b_0/comparator_0/AND_2/B Gnd 0.66fF
C4008 ALU_1b_0/AND_6/out Gnd 1.12fF
C4009 ALU_1b_0/comparator_0/AND_0/w_64_45# Gnd 1.05fF
C4010 ALU_1b_0/comparator_0/NOR_3/out Gnd 0.11fF
C4011 ALU_1b_0/comparator_0/NOR_3/A Gnd 1.06fF
C4012 ALU_1b_0/comparator_0/w_n195_n67# Gnd 1.09fF
C4013 ALU_1b_0/comparator_0/NOR_2/out Gnd 0.40fF
C4014 ALU_1b_0/comparator_0/NOR_2/B Gnd 1.06fF
C4015 ALU_1b_0/comparator_0/w_n220_n67# Gnd 1.09fF
C4016 ALU_1b_0/NOR_3/A Gnd 0.53fF
C4017 ALU_1b_0/AND_18/a_78_51# Gnd 0.42fF
C4018 ALU_1b_0/AND_18/w_64_45# Gnd 1.05fF
C4019 ALU_1b_0/NOR_0/A Gnd 0.80fF
C4020 ALU_1b_0/AND_19/a_78_51# Gnd 0.42fF
C4021 ALU_1b_0/AND_19/A Gnd 0.62fF
C4022 ALU_1b_0/AND_19/w_64_45# Gnd 1.05fF
C4023 ALU_1b_0/NOR_3/B Gnd 0.66fF
C4024 ALU_1b_0/AND_17/a_78_51# Gnd 0.42fF
C4025 ALU_1b_0/AND_17/w_64_45# Gnd 1.05fF
C4026 ALU_1b_0/NOR_0/B Gnd 0.69fF
C4027 ALU_1b_0/AND_16/a_78_51# Gnd 0.42fF
C4028 ALU_1b_0/AND_16/w_64_45# Gnd 1.05fF
C4029 ALU_1b_0/NOR_1/B Gnd 0.58fF
C4030 ALU_1b_0/AND_15/a_78_51# Gnd 0.42fF
C4031 ALU_1b_0/AND_15/w_64_45# Gnd 1.05fF
C4032 ALU_1b_0/AND_15/B Gnd 0.79fF
C4033 ALU_1b_0/AND_14/a_78_51# Gnd 0.42fF
C4034 ALU_1b_0/AND_14/B Gnd 0.93fF
C4035 ALU_1b_0/AND_14/A Gnd 0.42fF
C4036 ALU_1b_0/AND_9/a_78_51# Gnd 0.42fF
C4037 C1 Gnd 0.88fF
C4038 ALU_1b_0/AND_13/a_78_51# Gnd 0.42fF
C4039 ALU_1b_0/AND_14/w_64_45# Gnd 2.10fF
C4040 ALU_1b_0/AND_8/a_78_51# Gnd 0.42fF
C4041 C0 Gnd 0.95fF
C4042 ALU_1b_0/AND_8/w_64_45# Gnd 1.05fF
C4043 ALU_1b_0/AND_12/a_78_51# Gnd 0.42fF
C4044 ALU_1b_0/AND_7/a_78_51# Gnd 0.42fF
C4045 ALU_1b_0/AND_7/w_64_45# Gnd 1.05fF
C4046 ALU_1b_0/AND_6/a_78_51# Gnd 0.42fF
C4047 ALU_1b_0/AND_11/a_78_51# Gnd 0.42fF
C4048 ALU_1b_0/AND_10/a_78_51# Gnd 0.42fF
C4049 ALU_1b_0/AND_9/w_64_45# Gnd 3.15fF
C4050 ALU_1b_0/AND_4/a_78_51# Gnd 0.42fF
C4051 ALU_1b_0/AND_4/w_64_45# Gnd 1.05fF
C4052 ALU_1b_0/AND_5/a_78_51# Gnd 0.42fF
C4053 ALU_1b_0/AND_5/w_64_45# Gnd 1.05fF
C4054 ALU_1b_0/AND_3/a_78_51# Gnd 0.42fF
C4055 ALU_1b_0/AND_3/w_64_45# Gnd 1.53fF
C4056 ALU_1b_0/AND_2/a_78_51# Gnd 0.42fF
C4057 ALU_1b_0/AND_2/w_64_45# Gnd 1.05fF
C4058 ALU_1b_0/AND_18/A Gnd 0.73fF
C4059 ALU_1b_0/full_adder_1/NOR_0/out Gnd 0.39fF
C4060 ALU_1b_0/full_adder_1/w_448_45# Gnd 1.07fF
C4061 ALU_1b_0/full_adder_1/NOR_0/B Gnd 0.74fF
C4062 ALU_1b_0/AND_4/out Gnd 1.58fF
C4063 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C4064 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C4065 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C4066 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C4067 ALU_1b_0/AND_3/out Gnd 2.67fF
C4068 ALU_1b_0/full_adder_1/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C4069 ALU_1b_0/full_adder_1/half_adder_0/NAND_0/out Gnd 0.43fF
C4070 ALU_1b_0/full_adder_1/half_adder_0/w_36_45# Gnd 1.11fF
C4071 ALU_1b_0/full_adder_1/NOR_0/A Gnd 0.64fF
C4072 ALU_1b_0/AND_5/out Gnd 2.18fF
C4073 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C4074 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C4075 ALU_1b_0/NOT_1/in Gnd 1.41fF
C4076 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C4077 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C4078 ALU_1b_0/full_adder_1/half_adder_1/A Gnd 2.66fF
C4079 ALU_1b_0/full_adder_1/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C4080 ALU_1b_0/full_adder_1/half_adder_1/NAND_0/out Gnd 0.43fF
C4081 ALU_1b_0/full_adder_1/half_adder_1/w_36_45# Gnd 1.11fF
C4082 ALU_1b_0/AND_1/a_78_51# Gnd 0.42fF
C4083 ALU_1b_0/AND_1/w_64_45# Gnd 1.05fF
C4084 ALU_1b_0/AND_17/A Gnd 0.81fF
C4085 ALU_1b_0/full_adder_0/NOR_0/out Gnd 0.39fF
C4086 ALU_1b_0/full_adder_0/w_448_45# Gnd 1.07fF
C4087 ALU_1b_0/full_adder_0/NOR_0/B Gnd 0.74fF
C4088 ALU_1b_0/AND_2/out Gnd 1.53fF
C4089 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_177_36# Gnd 0.01fF
C4090 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_141_36# Gnd 0.01fF
C4091 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_184_44# Gnd 0.34fF
C4092 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/a_123_36# Gnd 0.80fF
C4093 ALU_1b_0/AND_0/out Gnd 3.03fF
C4094 ALU_1b_0/full_adder_0/half_adder_0/XOR_0/w_108_68# Gnd 2.10fF
C4095 ALU_1b_0/full_adder_0/half_adder_0/NAND_0/out Gnd 0.43fF
C4096 ALU_1b_0/full_adder_0/half_adder_0/w_36_45# Gnd 1.11fF
C4097 ALU_1b_0/full_adder_0/NOR_0/A Gnd 0.64fF
C4098 ALU_1b_0/AND_1/out Gnd 2.07fF
C4099 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_177_36# Gnd 0.01fF
C4100 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_141_36# Gnd 0.01fF
C4101 ALU_1b_0/AND_16/A Gnd 1.26fF
C4102 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_184_44# Gnd 0.34fF
C4103 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/a_123_36# Gnd 0.80fF
C4104 ALU_1b_0/full_adder_0/half_adder_1/A Gnd 2.66fF
C4105 ALU_1b_0/full_adder_0/half_adder_1/XOR_0/w_108_68# Gnd 2.10fF
C4106 ALU_1b_0/full_adder_0/half_adder_1/NAND_0/out Gnd 0.43fF
C4107 ALU_1b_0/full_adder_0/half_adder_1/w_36_45# Gnd 1.11fF
C4108 ALU_1b_0/AND_0/a_78_51# Gnd 0.42fF
C4109 ALU_1b_0/AND_0/w_64_45# Gnd 1.05fF
C4110 ALU_1b_0/NOT_6/in Gnd 0.42fF
C4111 ALU_1b_0/NOR_4/B Gnd 0.40fF
C4112 ALU_1b_0/NOR_4/A Gnd 0.82fF
C4113 ALU_1b_0/NOT_5/in Gnd 0.42fF
C4114 ALU_1b_0/NOR_4/w_n27_1# Gnd 2.18fF

***For Delay Analysis***

***For Subtraction wrt Cin***
Vin1 S0 GND supply
Vin2 S1 GND 0
Vin3 A0 GND 0
Vin4 A1 GND 0
Vin5 A2 GND 0
Vin6 A3 GND 0
Vin7 B0 GND 0
Vin8 B1 GND 0
Vin9 B2 GND 0
Vin10 B3 GND 0
Vin11 Cin GND pulse(0 supply 0 0.5p 0.5p 0.1u 0.2u)
Vin12 C1 GND 0
Vin13 C0 GND 0

.tran 1n 0.4u

.control
setplot const
run
echo "Delay due to Cin" > delay_analysis_sub_wrt_Cin.txt
meas tran trise00 trig v(Cin) val=0.5*supply rise=1 targ v(F0) val=0.5*supply rise=1
meas tran tfall00 trig v(Cin) val=0.5*supply fall=1 targ v(F0) val=0.5*supply fall=2
let tpd00 = (trise00 + tfall00)/2
echo "tpd00 = $&tpd00" >> delay_analysis_sub_wrt_Cin.txt
meas tran trise01 trig v(Cin) val=0.5*supply rise=1 targ v(F1) val=0.5*supply rise=1
meas tran tfall01 trig v(Cin) val=0.5*supply fall=1 targ v(F1) val=0.5*supply fall=2
let tpd01 = (trise01 + tfall01)/2
echo "tpd01 = $&tpd01" >> delay_analysis_sub_wrt_Cin.txt
meas tran trise02 trig v(Cin) val=0.5*supply rise=1 targ v(F2) val=0.5*supply rise=1
meas tran tfall02 trig v(Cin) val=0.5*supply fall=1 targ v(F2) val=0.5*supply fall=2
let tpd02 = (trise02 + tfall02)/2
echo "tpd02 = $&tpd02" >> delay_analysis_sub_wrt_Cin.txt
meas tran trise03 trig v(Cin) val=0.5*supply rise=1 targ v(F3) val=0.5*supply rise=1
meas tran tfall03 trig v(Cin) val=0.5*supply fall=1 targ v(F3) val=0.5*supply fall=2
let tpd03 = (trise03 + tfall03)/2
echo "tpd03 = $&tpd03" >> delay_analysis_sub_wrt_Cin.txt
meas tran trise04 trig v(Cin) val=0.5*supply rise=1 targ v(Cout) val=0.5*supply rise=1
meas tran tfall04 trig v(Cin) val=0.5*supply fall=1 targ v(Cout) val=0.5*supply fall=2
let tpd04 = (trise04 + tfall04)/2
echo "tpd04 = $&tpd04" >> delay_analysis_sub_wrt_Cin.txt
.endc

.end