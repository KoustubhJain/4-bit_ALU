*Two input CMOS NOR gate

.include TSMC_180nm.txt
.param supply=1.5
.option scale=0.09u

V1 vdd gnd supply

M1000 out B a_n14_10# vdd CMOSP w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1001 a_n14_10# A vdd vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1002 out A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=48 ps=40
M1003 gnd B out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A vdd 0.06fF
C1 A B 0.36fF
C2 A gnd 0.02fF
C3 vdd out 0.05fF
C4 vdd vdd 0.06fF
C5 vdd out 0.04fF
C6 out B 0.15fF
C7 vdd B 0.06fF
C8 gnd out 0.12fF
C9 gnd Gnd 0.16fF
C10 out Gnd 0.11fF
C11 vdd Gnd 0.05fF
C12 B Gnd 0.22fF
C13 A Gnd 0.21fF
C14 vdd Gnd 0.51fF

Vin1 A GND pulse(0 supply 0 0.5p 0.5p 0.1u 0.2u)
Vin2 B GND pulse(0 supply 0.15u 0.5p 0.5p 0.1u 0.2u)

.control
tran 1p 0.4u
plot v(A) v(B)+3 V(out)+6
.endc
.end