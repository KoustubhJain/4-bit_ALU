*Two input CMOS XOR gate

.include TSMC_180nm.txt
.param supply=1.5
.option scale=0.09u

V1 vdd gnd supply

M1000 out A a_141_36# Gnd CMOSN w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1001 a_123_36# A vdd vdd CMOSP w=4 l=2
+  ad=24 pd=20 as=104 ps=84
M1002 out B a_141_74# vdd CMOSP w=4 l=2
+  ad=44 pd=38 as=36 ps=26
M1003 a_141_36# B gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=104 ps=84
M1004 gnd a_184_44# a_177_36# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1005 a_141_74# a_123_36# vdd vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 vdd a_184_44# a_177_74# vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1007 a_177_36# a_123_36# out Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_177_74# A out vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 gnd B a_184_44# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1010 vdd B a_184_44# vdd CMOSP w=4 l=2
+  ad=0 pd=0 as=24 ps=20
M1011 a_123_36# A gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=0 ps=0
C0 out a_184_44# 0.13fF
C1 gnd A 0.03fF
C2 a_177_74# vdd 0.01fF
C3 out B 0.11fF
C4 vdd a_123_36# 0.06fF
C5 vdd vdd 0.23fF
C6 A a_123_36# 0.26fF
C7 B a_184_44# 0.06fF
C8 vdd A 0.13fF
C9 gnd a_141_36# 0.02fF
C10 gnd a_177_36# 0.02fF
C11 a_141_74# out 0.03fF
C12 vdd a_177_74# 0.02fF
C13 gnd a_184_44# 0.11fF
C14 out vdd 0.06fF
C15 vdd a_184_44# 0.09fF
C16 B a_123_36# 0.09fF
C17 vdd B 0.48fF
C18 out a_177_74# 0.03fF
C19 a_141_36# A 0.03fF
C20 gnd a_123_36# 0.14fF
C21 vdd a_184_44# 0.06fF
C22 out A 0.23fF
C23 a_141_74# vdd 0.01fF
C24 vdd B 0.06fF
C25 A a_184_44# 0.00fF
C26 vdd a_123_36# 0.09fF
C27 B A 0.08fF
C28 out a_141_36# 0.03fF
C29 out a_177_36# 0.03fF
C30 vdd a_141_74# 0.02fF
C31 a_177_36# Gnd 0.01fF
C32 a_141_36# Gnd 0.01fF
C33 gnd Gnd 0.25fF
C34 out Gnd 0.32fF
C35 vdd Gnd 0.10fF
C36 a_184_44# Gnd 0.34fF
C37 a_123_36# Gnd 0.80fF
C38 A Gnd 0.88fF
C39 B Gnd 0.26fF
C40 vdd Gnd 2.10fF

Vin1 A GND pulse(0 supply 0 0.5p 0.5p 0.1u 0.2u)
Vin2 B GND pulse(0 supply 0.15u 0.5p 0.5p 0.1u 0.2u)

.control
tran 1p 0.4u
plot v(A) v(B)+3 V(out)+6
.endc
.end