magic
tech scmos
timestamp 1701174042
<< nwell >>
rect -27 1 5 20
<< ntransistor >>
rect -16 -31 -14 -27
rect -8 -31 -6 -27
<< ptransistor >>
rect -16 7 -14 11
rect -8 7 -6 11
<< ndiffusion >>
rect -18 -31 -16 -27
rect -14 -31 -13 -27
rect -9 -31 -8 -27
rect -6 -31 -4 -27
<< pdiffusion >>
rect -17 7 -16 11
rect -14 7 -8 11
rect -6 7 -5 11
<< ndcontact >>
rect -22 -31 -18 -27
rect -13 -31 -9 -27
rect -4 -31 0 -27
<< pdcontact >>
rect -21 7 -17 11
rect -5 7 -1 11
<< polysilicon >>
rect -16 11 -14 14
rect -8 11 -6 14
rect -16 -27 -14 7
rect -8 -1 -6 7
rect -8 -27 -6 -5
rect -16 -34 -14 -31
rect -8 -34 -6 -31
<< polycontact >>
rect -20 -14 -16 -10
rect -10 -5 -6 -1
<< metal1 >>
rect -27 20 5 23
rect -21 11 -17 20
rect -1 -1 3 11
rect -27 -5 -10 -1
rect -1 -4 5 -1
rect -27 -14 -20 -10
rect -1 -12 3 -4
rect -13 -16 3 -12
rect -13 -27 -9 -16
rect -22 -40 -18 -31
rect -4 -40 0 -31
rect -27 -44 5 -40
<< labels >>
rlabel metal1 -19 21 -17 22 5 vdd
rlabel metal1 -25 -4 -23 -3 3 B
rlabel metal1 1 -3 3 -2 7 out
rlabel metal1 -12 -43 -10 -42 1 gnd
rlabel metal1 -26 -13 -24 -12 3 A
<< end >>
