CMOS Inverter
*Title

.include TSMC_180nm.txt
.param supply = 1.5
.option scale=0.09u
***Netlist***

Vdd vdd GND supply

M1000 out in vdd vdd CMOSP w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1001 out in gnd Gnd CMOSN w=4 l=2
+  ad=24 pd=20 as=20 ps=18
C0 in out 0.03fF
C1 vdd vdd 0.06fF
C2 out vdd 0.03fF
C3 gnd out 0.07fF
C4 out vdd 0.03fF
C5 in vdd 0.06fF
C6 gnd Gnd 0.06fF
C7 out Gnd 0.11fF
C8 vdd Gnd 0.02fF
C9 in Gnd 0.28fF
C10 vdd Gnd 0.48fF

Vin in GND pulse(0 supply 0 0.5p 0.5p 0.1u 0.2u)

.control
tran 1p 0.4u
plot v(out)+3 v(in)
.endc

.end
