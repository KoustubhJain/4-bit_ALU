magic
tech scmos
timestamp 1701520328
<< metal1 >>
rect 739 947 2162 951
rect 739 473 743 947
rect 1329 524 1333 947
rect 1356 876 1361 893
rect 1291 504 1421 509
rect 1291 415 1410 420
rect 149 220 158 224
rect 149 210 159 214
rect 149 196 158 200
rect 149 188 158 192
rect 149 180 159 184
rect 149 172 158 176
rect 1405 167 1410 415
rect 1416 185 1421 504
rect 2158 473 2162 947
rect 2711 504 2728 509
rect 2711 315 2716 420
rect 2615 310 2716 315
rect 1569 196 1579 200
rect 1569 188 1574 192
rect 1416 180 1574 185
rect 1552 177 1557 180
rect 1552 172 1575 177
rect 149 163 158 167
rect 1405 162 1575 167
rect 347 -169 350 23
rect 1329 -87 1333 -78
rect 1327 -91 1333 -87
rect 1327 -155 1331 -91
rect 1636 -166 1639 23
rect 1079 -169 1679 -166
rect 2615 -250 2620 310
rect 2723 304 2728 504
rect 1141 -255 1425 -250
rect 2561 -255 2620 -250
rect 2627 299 2728 304
rect 1141 -264 1415 -259
rect 1141 -272 1146 -264
rect 1141 -280 1145 -276
rect 1137 -288 1145 -284
rect -6 -508 -1 -503
rect -6 -597 -1 -592
rect 552 -991 556 -561
rect 1327 -991 1331 -276
rect 1410 -592 1415 -264
rect 1420 -508 1425 -255
rect 2627 -260 2632 299
rect 2562 -265 2632 -260
rect 2562 -272 2567 -265
rect 2558 -280 2566 -276
rect 2558 -288 2566 -284
rect 1410 -597 1425 -592
rect 1977 -991 1981 -565
rect 552 -995 1981 -991
<< m2contact >>
rect 1356 893 1361 898
rect 1356 871 1361 876
rect 1328 518 1334 524
rect 160 276 165 281
rect 168 265 173 270
rect 1580 289 1585 294
rect 1588 278 1593 283
rect 1328 -78 1334 -72
rect 1326 -161 1332 -155
rect 1326 -276 1332 -270
rect 1122 -339 1127 -334
rect 1130 -373 1135 -368
rect 2551 -328 2556 -323
rect 2543 -344 2548 -339
rect 2551 -370 2556 -365
rect 2543 -381 2548 -376
<< metal2 >>
rect -32 893 1356 898
rect 1361 893 2791 898
rect -32 270 -27 893
rect -17 882 2772 887
rect -17 281 -12 882
rect -17 276 160 281
rect -32 265 168 270
rect 1328 -72 1334 518
rect 1356 283 1361 871
rect 1393 294 1398 882
rect 1393 289 1580 294
rect 2767 283 2772 882
rect 1356 278 1588 283
rect 2667 278 2772 283
rect 1326 -270 1332 -161
rect 2667 -323 2672 278
rect 2786 258 2791 893
rect 2556 -328 2672 -323
rect 2691 253 2791 258
rect 1127 -339 1370 -334
rect 2691 -339 2696 253
rect 1135 -373 1331 -368
rect 1326 -959 1331 -373
rect 1365 -943 1370 -339
rect 2548 -344 2696 -339
rect 2556 -370 2737 -365
rect 2548 -381 2724 -376
rect 2719 -702 2724 -381
rect 2732 -686 2737 -370
rect 2732 -691 2754 -686
rect 2719 -707 2735 -702
rect 2730 -943 2735 -707
rect 1365 -948 2735 -943
rect 2749 -959 2754 -691
rect 1326 -964 2754 -959
use ALU_1b  ALU_1b_1
timestamp 1701510016
transform -1 0 1090 0 -1 -289
box -205 -201 1091 646
use ALU_1b  ALU_1b_3
timestamp 1701510016
transform -1 0 2511 0 -1 -289
box -205 -201 1091 646
use ALU_1b  ALU_1b_2
timestamp 1701510016
transform 1 0 1625 0 1 201
box -205 -201 1091 646
use ALU_1b  ALU_1b_0
timestamp 1701510016
transform 1 0 205 0 1 201
box -205 -201 1091 646
<< labels >>
rlabel metal1 1329 -135 1329 -135 1 gnd
rlabel metal1 1317 -168 1317 -168 1 vdd
rlabel metal1 150 198 150 198 1 A0
rlabel metal1 150 190 150 190 1 B0
rlabel metal1 150 182 150 182 1 Cin
rlabel metal1 150 174 150 174 1 C0
rlabel metal1 150 165 150 165 1 C1
rlabel metal1 150 222 150 222 1 S1
rlabel metal1 150 212 150 212 1 S0
rlabel metal1 1305 417 1305 417 1 F0
rlabel metal1 1570 198 1570 198 1 A1
rlabel metal1 1570 190 1570 190 1 B1
rlabel metal1 2713 388 2713 388 1 F1
rlabel metal1 2564 -286 2564 -286 1 A2
rlabel metal1 2564 -278 2564 -278 1 B2
rlabel metal1 1422 -482 1422 -482 1 F2
rlabel metal1 1144 -286 1144 -286 1 A3
rlabel metal1 1144 -278 1144 -278 1 B3
rlabel metal1 -5 -505 -5 -505 1 F3
rlabel metal1 -5 -594 -5 -594 1 Cout
<< end >>
